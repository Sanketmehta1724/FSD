<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>2.69797,-144.53,91.9698,-188.656</PageViewport>
<gate>
<ID>2</ID>
<type>BA_NAND2</type>
<position>30,-13</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>BA_NAND2</type>
<position>29.5,-23</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>BA_NAND2</type>
<position>51,-13</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8</ID>
<type>BA_NAND2</type>
<position>51,-22</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>14.5,-7</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>12</ID>
<type>GA_LED</type>
<position>63,-13</position>
<input>
<ID>N_in0</ID>4 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>GA_LED</type>
<position>63.5,-22</position>
<input>
<ID>N_in0</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>BB_CLOCK</type>
<position>20,-18</position>
<output>
<ID>CLK</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 60</lparam></gate>
<gate>
<ID>20</ID>
<type>AE_SMALL_INVERTER</type>
<position>14.5,-12.5</position>
<input>
<ID>IN_0</ID>6 </input>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>23</ID>
<type>AA_TOGGLE</type>
<position>80.5,-12.5</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>24</ID>
<type>BB_CLOCK</type>
<position>82,-17.5</position>
<output>
<ID>CLK</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 60</lparam></gate>
<gate>
<ID>26</ID>
<type>GA_LED</type>
<position>100,-14</position>
<input>
<ID>N_in0</ID>16 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>219</ID>
<type>AA_LABEL</type>
<position>-13.5,-153</position>
<gparam>LABEL_TEXT SR TO JKFF</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>27</ID>
<type>GA_LED</type>
<position>100.5,-23</position>
<input>
<ID>N_in0</ID>15 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>29</ID>
<type>AE_DFF_LOW</type>
<position>91,-16.5</position>
<input>
<ID>IN_0</ID>13 </input>
<output>
<ID>OUTINV_0</ID>15 </output>
<output>
<ID>OUT_0</ID>16 </output>
<input>
<ID>clock</ID>14 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>31</ID>
<type>AA_LABEL</type>
<position>60.5,-4.5</position>
<gparam>LABEL_TEXT D FF</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>AA_LABEL</type>
<position>15,-4.5</position>
<gparam>LABEL_TEXT D </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>33</ID>
<type>AA_LABEL</type>
<position>66.5,-13</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>34</ID>
<type>AA_LABEL</type>
<position>67,-21.5</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>AA_LABEL</type>
<position>67,-18.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>AA_LABEL</type>
<position>105,-13.5</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>37</ID>
<type>AA_LABEL</type>
<position>105.5,-22</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>AA_LABEL</type>
<position>105.5,-19</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>AA_LABEL</type>
<position>77.5,-12</position>
<gparam>LABEL_TEXT D </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>41</ID>
<type>BE_JKFF_LOW</type>
<position>25,-37</position>
<input>
<ID>J</ID>18 </input>
<input>
<ID>K</ID>19 </input>
<output>
<ID>Q</ID>20 </output>
<input>
<ID>clock</ID>17 </input>
<output>
<ID>nQ</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>43</ID>
<type>AA_TOGGLE</type>
<position>11.5,-33.5</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>45</ID>
<type>AA_TOGGLE</type>
<position>11,-40</position>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>47</ID>
<type>BB_CLOCK</type>
<position>16.5,-37</position>
<output>
<ID>CLK</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 60</lparam></gate>
<gate>
<ID>50</ID>
<type>GA_LED</type>
<position>35,-33</position>
<input>
<ID>N_in0</ID>20 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>51</ID>
<type>GA_LED</type>
<position>35.5,-42</position>
<input>
<ID>N_in0</ID>21 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>52</ID>
<type>AA_LABEL</type>
<position>40,-32.5</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>53</ID>
<type>AA_LABEL</type>
<position>40.5,-41</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>54</ID>
<type>AA_LABEL</type>
<position>40.5,-38</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>55</ID>
<type>AA_LABEL</type>
<position>23.5,-28.5</position>
<gparam>LABEL_TEXT JK FF</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>56</ID>
<type>AA_LABEL</type>
<position>8,-33</position>
<gparam>LABEL_TEXT J</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>57</ID>
<type>AA_LABEL</type>
<position>7.5,-39.5</position>
<gparam>LABEL_TEXT K</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>58</ID>
<type>BE_JKFF_LOW</type>
<position>92.5,-38</position>
<input>
<ID>J</ID>23 </input>
<input>
<ID>K</ID>23 </input>
<output>
<ID>Q</ID>25 </output>
<input>
<ID>clock</ID>22 </input>
<output>
<ID>nQ</ID>26 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>59</ID>
<type>AA_TOGGLE</type>
<position>77.5,-32</position>
<output>
<ID>OUT_0</ID>23 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>61</ID>
<type>BB_CLOCK</type>
<position>84,-38</position>
<output>
<ID>CLK</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 60</lparam></gate>
<gate>
<ID>62</ID>
<type>GA_LED</type>
<position>102.5,-34</position>
<input>
<ID>N_in0</ID>25 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>63</ID>
<type>GA_LED</type>
<position>103,-43</position>
<input>
<ID>N_in0</ID>26 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>64</ID>
<type>AA_LABEL</type>
<position>107.5,-33.5</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>65</ID>
<type>AA_LABEL</type>
<position>108,-42</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>66</ID>
<type>AA_LABEL</type>
<position>108,-39</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>67</ID>
<type>AA_LABEL</type>
<position>74.5,-31.5</position>
<gparam>LABEL_TEXT T</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>69</ID>
<type>AA_LABEL</type>
<position>87.5,-27.5</position>
<gparam>LABEL_TEXT T FF</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>AA_LABEL</type>
<position>20.5,-48.5</position>
<gparam>LABEL_TEXT D TO SR FF</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>71</ID>
<type>AA_TOGGLE</type>
<position>-10.5,-53</position>
<output>
<ID>OUT_0</ID>34 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>72</ID>
<type>BB_CLOCK</type>
<position>8.5,-60.5</position>
<output>
<ID>CLK</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 60</lparam></gate>
<gate>
<ID>73</ID>
<type>GA_LED</type>
<position>26.5,-57</position>
<input>
<ID>N_in0</ID>30 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>74</ID>
<type>GA_LED</type>
<position>27,-66</position>
<input>
<ID>N_in0</ID>29 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>75</ID>
<type>AE_DFF_LOW</type>
<position>17.5,-59.5</position>
<input>
<ID>IN_0</ID>36 </input>
<output>
<ID>OUTINV_0</ID>29 </output>
<output>
<ID>OUT_0</ID>30 </output>
<input>
<ID>clock</ID>28 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>76</ID>
<type>AA_LABEL</type>
<position>31.5,-56.5</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>77</ID>
<type>AA_LABEL</type>
<position>32,-65</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>78</ID>
<type>AA_LABEL</type>
<position>32,-62</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>81</ID>
<type>AA_AND2</type>
<position>-3.5,-59</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>30 </input>
<output>
<ID>OUT</ID>35 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>83</ID>
<type>AE_OR2</type>
<position>8,-54.5</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>35 </input>
<output>
<ID>OUT</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>85</ID>
<type>AA_TOGGLE</type>
<position>-15,-58</position>
<output>
<ID>OUT_0</ID>33 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>87</ID>
<type>AE_SMALL_INVERTER</type>
<position>-10,-58</position>
<input>
<ID>IN_0</ID>33 </input>
<output>
<ID>OUT_0</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>97</ID>
<type>AA_LABEL</type>
<position>92,-48.5</position>
<gparam>LABEL_TEXT D TO JK FF</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>98</ID>
<type>AA_TOGGLE</type>
<position>67.5,-56</position>
<output>
<ID>OUT_0</ID>49 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>99</ID>
<type>BB_CLOCK</type>
<position>91.5,-61.5</position>
<output>
<ID>CLK</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 60</lparam></gate>
<gate>
<ID>100</ID>
<type>GA_LED</type>
<position>109.5,-58</position>
<input>
<ID>N_in0</ID>43 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>101</ID>
<type>GA_LED</type>
<position>110,-67</position>
<input>
<ID>N_in0</ID>42 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>102</ID>
<type>AE_DFF_LOW</type>
<position>100.5,-60.5</position>
<input>
<ID>IN_0</ID>48 </input>
<output>
<ID>OUTINV_0</ID>42 </output>
<output>
<ID>OUT_0</ID>43 </output>
<input>
<ID>clock</ID>41 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 0</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>103</ID>
<type>AA_LABEL</type>
<position>114.5,-57.5</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>104</ID>
<type>AA_LABEL</type>
<position>115,-66</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>105</ID>
<type>AA_LABEL</type>
<position>115,-63</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>106</ID>
<type>AA_AND2</type>
<position>79.5,-60</position>
<input>
<ID>IN_0</ID>44 </input>
<input>
<ID>IN_1</ID>43 </input>
<output>
<ID>OUT</ID>47 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>107</ID>
<type>AE_OR2</type>
<position>91,-55.5</position>
<input>
<ID>IN_0</ID>50 </input>
<input>
<ID>IN_1</ID>47 </input>
<output>
<ID>OUT</ID>48 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>108</ID>
<type>AA_TOGGLE</type>
<position>68,-59</position>
<output>
<ID>OUT_0</ID>45 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>109</ID>
<type>AE_SMALL_INVERTER</type>
<position>73,-59</position>
<input>
<ID>IN_0</ID>45 </input>
<output>
<ID>OUT_0</ID>44 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>111</ID>
<type>AA_AND2</type>
<position>77,-55</position>
<input>
<ID>IN_0</ID>42 </input>
<input>
<ID>IN_1</ID>49 </input>
<output>
<ID>OUT</ID>50 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>112</ID>
<type>AA_LABEL</type>
<position>51.5,-73.5</position>
<gparam>LABEL_TEXT D TO T FF</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>114</ID>
<type>BB_CLOCK</type>
<position>51,-86.5</position>
<output>
<ID>CLK</ID>51 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 60</lparam></gate>
<gate>
<ID>115</ID>
<type>GA_LED</type>
<position>69,-83</position>
<input>
<ID>N_in0</ID>53 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>116</ID>
<type>GA_LED</type>
<position>69.5,-92</position>
<input>
<ID>N_in0</ID>52 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>117</ID>
<type>AE_DFF_LOW</type>
<position>60,-85.5</position>
<input>
<ID>IN_0</ID>61 </input>
<output>
<ID>OUTINV_0</ID>52 </output>
<output>
<ID>OUT_0</ID>53 </output>
<input>
<ID>clock</ID>51 </input>
<gparam>angle 0.0</gparam>
<lparam>CURRENT_VALUE 1</lparam>
<lparam>INPUT_BITS 1</lparam>
<lparam>NO_HOLD true</lparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_LOAD true</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>118</ID>
<type>AA_LABEL</type>
<position>74,-82.5</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>119</ID>
<type>AA_LABEL</type>
<position>74.5,-91</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>120</ID>
<type>AA_LABEL</type>
<position>74.5,-88</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>127</ID>
<type>AI_XOR2</type>
<position>48,-82</position>
<input>
<ID>IN_0</ID>53 </input>
<input>
<ID>IN_1</ID>60 </input>
<output>
<ID>OUT</ID>61 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>129</ID>
<type>AA_TOGGLE</type>
<position>37.5,-83</position>
<output>
<ID>OUT_0</ID>60 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>130</ID>
<type>BE_JKFF_LOW</type>
<position>-8.5,-105.5</position>
<input>
<ID>J</ID>63 </input>
<input>
<ID>K</ID>64 </input>
<output>
<ID>Q</ID>65 </output>
<input>
<ID>clock</ID>62 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>131</ID>
<type>AA_TOGGLE</type>
<position>-22,-102</position>
<output>
<ID>OUT_0</ID>63 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>132</ID>
<type>AA_TOGGLE</type>
<position>-22.5,-108.5</position>
<output>
<ID>OUT_0</ID>64 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>133</ID>
<type>BB_CLOCK</type>
<position>-17,-105.5</position>
<output>
<ID>CLK</ID>62 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 60</lparam></gate>
<gate>
<ID>134</ID>
<type>GA_LED</type>
<position>1.5,-101.5</position>
<input>
<ID>N_in0</ID>65 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>136</ID>
<type>AA_LABEL</type>
<position>6.5,-101</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>139</ID>
<type>AA_LABEL</type>
<position>-25.5,-101.5</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>140</ID>
<type>AA_LABEL</type>
<position>-26,-108</position>
<gparam>LABEL_TEXT R</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>141</ID>
<type>AA_LABEL</type>
<position>-11.5,-96</position>
<gparam>LABEL_TEXT JK TO SR FF</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>156</ID>
<type>BE_JKFF_LOW</type>
<position>39,-105.5</position>
<input>
<ID>J</ID>76 </input>
<input>
<ID>K</ID>80 </input>
<output>
<ID>Q</ID>78 </output>
<input>
<ID>clock</ID>75 </input>
<output>
<ID>nQ</ID>79 </output>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>157</ID>
<type>AA_TOGGLE</type>
<position>25,-101.5</position>
<output>
<ID>OUT_0</ID>76 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>159</ID>
<type>BB_CLOCK</type>
<position>29.5,-106</position>
<output>
<ID>CLK</ID>75 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 60</lparam></gate>
<gate>
<ID>160</ID>
<type>GA_LED</type>
<position>49,-101.5</position>
<input>
<ID>N_in0</ID>78 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>161</ID>
<type>AA_LABEL</type>
<position>54,-101</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>162</ID>
<type>AA_LABEL</type>
<position>38,-95</position>
<gparam>LABEL_TEXT JK TO D FF</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>163</ID>
<type>GA_LED</type>
<position>49,-107.5</position>
<input>
<ID>N_in0</ID>79 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>164</ID>
<type>AA_LABEL</type>
<position>54,-107</position>
<gparam>LABEL_TEXT Q'</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>166</ID>
<type>AE_OR2</type>
<position>26.5,-110</position>
<input>
<ID>IN_0</ID>76 </input>
<input>
<ID>IN_1</ID>79 </input>
<output>
<ID>OUT</ID>80 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>169</ID>
<type>BE_JKFF_LOW</type>
<position>-9.5,-136.5</position>
<input>
<ID>J</ID>85 </input>
<input>
<ID>K</ID>85 </input>
<output>
<ID>Q</ID>84 </output>
<input>
<ID>clock</ID>81 </input>
<gparam>angle 0.0</gparam>
<lparam>SYNC_CLEAR false</lparam>
<lparam>SYNC_SET false</lparam></gate>
<gate>
<ID>170</ID>
<type>AA_TOGGLE</type>
<position>-26,-132</position>
<output>
<ID>OUT_0</ID>85 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>172</ID>
<type>BB_CLOCK</type>
<position>-18,-136.5</position>
<output>
<ID>CLK</ID>81 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 60</lparam></gate>
<gate>
<ID>173</ID>
<type>GA_LED</type>
<position>0.5,-132.5</position>
<input>
<ID>N_in0</ID>84 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>174</ID>
<type>AA_LABEL</type>
<position>5.5,-132</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>175</ID>
<type>AA_LABEL</type>
<position>-26,-129</position>
<gparam>LABEL_TEXT T</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>177</ID>
<type>AA_LABEL</type>
<position>-12.5,-127</position>
<gparam>LABEL_TEXT JK TO T FF</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>178</ID>
<type>BA_NAND2</type>
<position>44,-132</position>
<input>
<ID>IN_0</ID>91 </input>
<input>
<ID>IN_1</ID>90 </input>
<output>
<ID>OUT</ID>86 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>179</ID>
<type>BA_NAND2</type>
<position>43.5,-142</position>
<input>
<ID>IN_0</ID>90 </input>
<input>
<ID>IN_1</ID>92 </input>
<output>
<ID>OUT</ID>87 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>180</ID>
<type>BA_NAND2</type>
<position>65,-132</position>
<input>
<ID>IN_0</ID>86 </input>
<input>
<ID>IN_1</ID>88 </input>
<output>
<ID>OUT</ID>89 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>181</ID>
<type>BA_NAND2</type>
<position>65,-141</position>
<input>
<ID>IN_0</ID>89 </input>
<input>
<ID>IN_1</ID>87 </input>
<output>
<ID>OUT</ID>88 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>182</ID>
<type>AA_TOGGLE</type>
<position>28.5,-126</position>
<output>
<ID>OUT_0</ID>91 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>183</ID>
<type>GA_LED</type>
<position>77,-132</position>
<input>
<ID>N_in0</ID>89 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>184</ID>
<type>GA_LED</type>
<position>77.5,-141</position>
<input>
<ID>N_in0</ID>88 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>185</ID>
<type>BB_CLOCK</type>
<position>34,-137</position>
<output>
<ID>CLK</ID>90 </output>
<gparam>angle 0.0</gparam>
<lparam>HALF_CYCLE 60</lparam></gate>
<gate>
<ID>186</ID>
<type>AE_SMALL_INVERTER</type>
<position>28.5,-131.5</position>
<input>
<ID>IN_0</ID>91 </input>
<output>
<ID>OUT_0</ID>92 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>187</ID>
<type>AA_LABEL</type>
<position>74.5,-123.5</position>
<gparam>LABEL_TEXT SR TO D FF</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>188</ID>
<type>AA_LABEL</type>
<position>29,-123.5</position>
<gparam>LABEL_TEXT D </gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>189</ID>
<type>AA_LABEL</type>
<position>80.5,-132</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>190</ID>
<type>AA_LABEL</type>
<position>81,-140.5</position>
<gparam>LABEL_TEXT Q</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>191</ID>
<type>AA_LABEL</type>
<position>81,-137.5</position>
<gparam>LABEL_TEXT _</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-13,40.5,-12</points>
<intersection>-13 2</intersection>
<intersection>-12 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,-12,48,-12</points>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>33,-13,40.5,-13</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<intersection>40.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>32.5,-23,48,-23</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<connection>
<GID>4</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54,-22,62.5,-22</points>
<connection>
<GID>8</GID>
<name>OUT</name></connection>
<connection>
<GID>14</GID>
<name>N_in0</name></connection>
<intersection>55 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>55,-22,55,-16.5</points>
<intersection>-22 1</intersection>
<intersection>-16.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>48,-16.5,55,-16.5</points>
<intersection>48 5</intersection>
<intersection>55 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>48,-16.5,48,-14</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>-16.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54,-13,62,-13</points>
<connection>
<GID>12</GID>
<name>N_in0</name></connection>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<intersection>54.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>54.5,-19,54.5,-13</points>
<intersection>-19 4</intersection>
<intersection>-13 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>48,-19,54.5,-19</points>
<intersection>48 5</intersection>
<intersection>54.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>48,-21,48,-19</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>-19 4</intersection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>26.5,-22,26.5,-14</points>
<connection>
<GID>4</GID>
<name>IN_0</name></connection>
<intersection>-18 2</intersection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>26.5,-14,27,-14</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<intersection>26.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>24,-18,26.5,-18</points>
<connection>
<GID>16</GID>
<name>CLK</name></connection>
<intersection>26.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-10.5,14.5,-9</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>-10 3</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>14.5,-10,27,-10</points>
<intersection>14.5 0</intersection>
<intersection>27 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>27,-12,27,-10</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>-10 3</intersection></vsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>14.5,-24,14.5,-14.5</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>-24 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>14.5,-24,26.5,-24</points>
<connection>
<GID>4</GID>
<name>IN_1</name></connection>
<intersection>14.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,-14.5,85,-12.5</points>
<intersection>-14.5 1</intersection>
<intersection>-12.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85,-14.5,88,-14.5</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<intersection>85 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>82.5,-12.5,85,-12.5</points>
<connection>
<GID>23</GID>
<name>OUT_0</name></connection>
<intersection>85 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>86,-17.5,88,-17.5</points>
<connection>
<GID>24</GID>
<name>CLK</name></connection>
<connection>
<GID>29</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96.5,-23,96.5,-17.5</points>
<intersection>-23 1</intersection>
<intersection>-17.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>96.5,-23,99.5,-23</points>
<connection>
<GID>27</GID>
<name>N_in0</name></connection>
<intersection>96.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>94,-17.5,96.5,-17.5</points>
<connection>
<GID>29</GID>
<name>OUTINV_0</name></connection>
<intersection>96.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>96.5,-14.5,96.5,-14</points>
<intersection>-14.5 2</intersection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>96.5,-14,99,-14</points>
<connection>
<GID>26</GID>
<name>N_in0</name></connection>
<intersection>96.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>94,-14.5,96.5,-14.5</points>
<connection>
<GID>29</GID>
<name>OUT_0</name></connection>
<intersection>96.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20.5,-37,22,-37</points>
<connection>
<GID>41</GID>
<name>clock</name></connection>
<connection>
<GID>47</GID>
<name>CLK</name></connection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13.5,-33.5,22,-33.5</points>
<connection>
<GID>43</GID>
<name>OUT_0</name></connection>
<intersection>22 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>22,-35,22,-33.5</points>
<connection>
<GID>41</GID>
<name>J</name></connection>
<intersection>-33.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>13,-40,22,-40</points>
<connection>
<GID>45</GID>
<name>OUT_0</name></connection>
<intersection>22 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>22,-40,22,-39</points>
<connection>
<GID>41</GID>
<name>K</name></connection>
<intersection>-40 1</intersection></vsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-35,31,-33</points>
<intersection>-35 2</intersection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-33,34,-33</points>
<connection>
<GID>50</GID>
<name>N_in0</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28,-35,31,-35</points>
<connection>
<GID>41</GID>
<name>Q</name></connection>
<intersection>31 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-42,31,-39</points>
<intersection>-42 1</intersection>
<intersection>-39 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-42,34.5,-42</points>
<connection>
<GID>51</GID>
<name>N_in0</name></connection>
<intersection>31 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>28,-39,31,-39</points>
<connection>
<GID>41</GID>
<name>nQ</name></connection>
<intersection>31 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>88,-38,89.5,-38</points>
<connection>
<GID>58</GID>
<name>clock</name></connection>
<connection>
<GID>61</GID>
<name>CLK</name></connection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>79.5,-32,80,-32</points>
<connection>
<GID>59</GID>
<name>OUT_0</name></connection>
<intersection>80 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>80,-40,80,-32</points>
<intersection>-40 5</intersection>
<intersection>-36 6</intersection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>80,-40,89.5,-40</points>
<connection>
<GID>58</GID>
<name>K</name></connection>
<intersection>80 3</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>80,-36,89.5,-36</points>
<connection>
<GID>58</GID>
<name>J</name></connection>
<intersection>80 3</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98.5,-36,98.5,-34</points>
<intersection>-36 2</intersection>
<intersection>-34 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98.5,-34,101.5,-34</points>
<connection>
<GID>62</GID>
<name>N_in0</name></connection>
<intersection>98.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>95.5,-36,98.5,-36</points>
<connection>
<GID>58</GID>
<name>Q</name></connection>
<intersection>98.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>98.5,-43,98.5,-40</points>
<intersection>-43 1</intersection>
<intersection>-40 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>98.5,-43,102,-43</points>
<connection>
<GID>63</GID>
<name>N_in0</name></connection>
<intersection>98.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>95.5,-40,98.5,-40</points>
<connection>
<GID>58</GID>
<name>nQ</name></connection>
<intersection>98.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>12.5,-60.5,14.5,-60.5</points>
<connection>
<GID>72</GID>
<name>CLK</name></connection>
<connection>
<GID>75</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>23,-66,23,-60.5</points>
<intersection>-66 1</intersection>
<intersection>-60.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>23,-66,26,-66</points>
<connection>
<GID>74</GID>
<name>N_in0</name></connection>
<intersection>23 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>20.5,-60.5,23,-60.5</points>
<connection>
<GID>75</GID>
<name>OUTINV_0</name></connection>
<intersection>23 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>20.5,-66,20.5,-57</points>
<connection>
<GID>75</GID>
<name>OUT_0</name></connection>
<intersection>-66 2</intersection>
<intersection>-57 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>20.5,-57,25.5,-57</points>
<connection>
<GID>73</GID>
<name>N_in0</name></connection>
<intersection>20.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-6.5,-66,20.5,-66</points>
<intersection>-6.5 3</intersection>
<intersection>20.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-6.5,-66,-6.5,-60</points>
<connection>
<GID>81</GID>
<name>IN_1</name></connection>
<intersection>-66 2</intersection></vsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-8,-58,-6.5,-58</points>
<connection>
<GID>87</GID>
<name>OUT_0</name></connection>
<connection>
<GID>81</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13,-58,-12,-58</points>
<connection>
<GID>85</GID>
<name>OUT_0</name></connection>
<connection>
<GID>87</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-1.5,-53.5,-1.5,-53</points>
<intersection>-53.5 1</intersection>
<intersection>-53 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-1.5,-53.5,5,-53.5</points>
<connection>
<GID>83</GID>
<name>IN_0</name></connection>
<intersection>-1.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-8.5,-53,-1.5,-53</points>
<connection>
<GID>71</GID>
<name>OUT_0</name></connection>
<intersection>-1.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>2,-59,2,-55.5</points>
<intersection>-59 2</intersection>
<intersection>-55.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>2,-55.5,5,-55.5</points>
<connection>
<GID>83</GID>
<name>IN_1</name></connection>
<intersection>2 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-0.5,-59,2,-59</points>
<connection>
<GID>81</GID>
<name>OUT</name></connection>
<intersection>2 0</intersection></hsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>12.5,-57.5,12.5,-54.5</points>
<intersection>-57.5 1</intersection>
<intersection>-54.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>12.5,-57.5,14.5,-57.5</points>
<connection>
<GID>75</GID>
<name>IN_0</name></connection>
<intersection>12.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>11,-54.5,12.5,-54.5</points>
<connection>
<GID>83</GID>
<name>OUT</name></connection>
<intersection>12.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>95.5,-61.5,97.5,-61.5</points>
<connection>
<GID>99</GID>
<name>CLK</name></connection>
<connection>
<GID>102</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106.5,-67,106.5,-51.5</points>
<intersection>-67 1</intersection>
<intersection>-61.5 5</intersection>
<intersection>-51.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>106.5,-67,109,-67</points>
<connection>
<GID>101</GID>
<name>N_in0</name></connection>
<intersection>106.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>74,-51.5,106.5,-51.5</points>
<intersection>74 3</intersection>
<intersection>106.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>74,-54,74,-51.5</points>
<connection>
<GID>111</GID>
<name>IN_0</name></connection>
<intersection>-51.5 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>103.5,-61.5,106.5,-61.5</points>
<connection>
<GID>102</GID>
<name>OUTINV_0</name></connection>
<intersection>106.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104,-67,104,-58</points>
<intersection>-67 2</intersection>
<intersection>-58.5 4</intersection>
<intersection>-58 5</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>76.5,-67,104,-67</points>
<intersection>76.5 3</intersection>
<intersection>104 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>76.5,-67,76.5,-61</points>
<connection>
<GID>106</GID>
<name>IN_1</name></connection>
<intersection>-67 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>103.5,-58.5,104,-58.5</points>
<connection>
<GID>102</GID>
<name>OUT_0</name></connection>
<intersection>104 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>104,-58,108.5,-58</points>
<connection>
<GID>100</GID>
<name>N_in0</name></connection>
<intersection>104 0</intersection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>75,-59,76.5,-59</points>
<connection>
<GID>109</GID>
<name>OUT_0</name></connection>
<connection>
<GID>106</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>70,-59,71,-59</points>
<connection>
<GID>108</GID>
<name>OUT_0</name></connection>
<connection>
<GID>109</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,-60,85,-56.5</points>
<intersection>-60 2</intersection>
<intersection>-56.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85,-56.5,88,-56.5</points>
<connection>
<GID>107</GID>
<name>IN_1</name></connection>
<intersection>85 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>82.5,-60,85,-60</points>
<connection>
<GID>106</GID>
<name>OUT</name></connection>
<intersection>85 0</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>95.5,-58.5,95.5,-55.5</points>
<intersection>-58.5 1</intersection>
<intersection>-55.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>95.5,-58.5,97.5,-58.5</points>
<connection>
<GID>102</GID>
<name>IN_0</name></connection>
<intersection>95.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>94,-55.5,95.5,-55.5</points>
<connection>
<GID>107</GID>
<name>OUT</name></connection>
<intersection>95.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>69.5,-56,74,-56</points>
<connection>
<GID>98</GID>
<name>OUT_0</name></connection>
<connection>
<GID>111</GID>
<name>IN_1</name></connection></hsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>84,-55,84,-54.5</points>
<intersection>-55 2</intersection>
<intersection>-54.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>84,-54.5,88,-54.5</points>
<connection>
<GID>107</GID>
<name>IN_0</name></connection>
<intersection>84 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>80,-55,84,-55</points>
<connection>
<GID>111</GID>
<name>OUT</name></connection>
<intersection>84 0</intersection></hsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>55,-86.5,57,-86.5</points>
<connection>
<GID>117</GID>
<name>clock</name></connection>
<connection>
<GID>114</GID>
<name>CLK</name></connection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66,-92,66,-86.5</points>
<intersection>-92 1</intersection>
<intersection>-86.5 5</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66,-92,68.5,-92</points>
<connection>
<GID>116</GID>
<name>N_in0</name></connection>
<intersection>66 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>63,-86.5,66,-86.5</points>
<connection>
<GID>117</GID>
<name>OUTINV_0</name></connection>
<intersection>66 0</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>63.5,-83.5,63.5,-79</points>
<intersection>-83.5 9</intersection>
<intersection>-83 5</intersection>
<intersection>-79 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>45,-79,63.5,-79</points>
<intersection>45 7</intersection>
<intersection>63.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>63.5,-83,68,-83</points>
<connection>
<GID>115</GID>
<name>N_in0</name></connection>
<intersection>63.5 0</intersection></hsegment>
<vsegment>
<ID>7</ID>
<points>45,-81,45,-79</points>
<connection>
<GID>127</GID>
<name>IN_0</name></connection>
<intersection>-79 4</intersection></vsegment>
<hsegment>
<ID>9</ID>
<points>63,-83.5,63.5,-83.5</points>
<connection>
<GID>117</GID>
<name>OUT_0</name></connection>
<intersection>63.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39.5,-83,45,-83</points>
<connection>
<GID>127</GID>
<name>IN_1</name></connection>
<connection>
<GID>129</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-83.5,54,-82</points>
<intersection>-83.5 1</intersection>
<intersection>-82 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54,-83.5,57,-83.5</points>
<connection>
<GID>117</GID>
<name>IN_0</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>51,-82,54,-82</points>
<connection>
<GID>127</GID>
<name>OUT</name></connection>
<intersection>54 0</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-13,-105.5,-11.5,-105.5</points>
<connection>
<GID>133</GID>
<name>CLK</name></connection>
<connection>
<GID>130</GID>
<name>clock</name></connection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-20,-102,-11.5,-102</points>
<connection>
<GID>131</GID>
<name>OUT_0</name></connection>
<intersection>-11.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-11.5,-103.5,-11.5,-102</points>
<connection>
<GID>130</GID>
<name>J</name></connection>
<intersection>-102 1</intersection></vsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-20.5,-108.5,-11.5,-108.5</points>
<connection>
<GID>132</GID>
<name>OUT_0</name></connection>
<intersection>-11.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-11.5,-108.5,-11.5,-107.5</points>
<connection>
<GID>130</GID>
<name>K</name></connection>
<intersection>-108.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-2.5,-103.5,-2.5,-101.5</points>
<intersection>-103.5 2</intersection>
<intersection>-101.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-2.5,-101.5,0.5,-101.5</points>
<connection>
<GID>134</GID>
<name>N_in0</name></connection>
<intersection>-2.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-5.5,-103.5,-2.5,-103.5</points>
<connection>
<GID>130</GID>
<name>Q</name></connection>
<intersection>-2.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>33.5,-106,36,-106</points>
<connection>
<GID>159</GID>
<name>CLK</name></connection>
<intersection>36 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>36,-106,36,-105.5</points>
<connection>
<GID>156</GID>
<name>clock</name></connection>
<intersection>-106 1</intersection></vsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>20,-100,28,-100</points>
<intersection>20 4</intersection>
<intersection>28 6</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>20,-109,20,-100</points>
<intersection>-109 10</intersection>
<intersection>-100 1</intersection></vsegment>
<vsegment>
<ID>6</ID>
<points>28,-103.5,28,-100</points>
<intersection>-103.5 9</intersection>
<intersection>-101.5 8</intersection>
<intersection>-100 1</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>27,-101.5,28,-101.5</points>
<connection>
<GID>157</GID>
<name>OUT_0</name></connection>
<intersection>28 6</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>28,-103.5,36,-103.5</points>
<connection>
<GID>156</GID>
<name>J</name></connection>
<intersection>28 6</intersection></hsegment>
<hsegment>
<ID>10</ID>
<points>20,-109,23.5,-109</points>
<connection>
<GID>166</GID>
<name>IN_0</name></connection>
<intersection>20 4</intersection></hsegment></shape></wire>
<wire>
<ID>78</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>45,-103.5,45,-101.5</points>
<intersection>-103.5 2</intersection>
<intersection>-101.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>45,-101.5,48,-101.5</points>
<connection>
<GID>160</GID>
<name>N_in0</name></connection>
<intersection>45 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>42,-103.5,45,-103.5</points>
<connection>
<GID>156</GID>
<name>Q</name></connection>
<intersection>45 0</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>23.5,-111,48,-111</points>
<connection>
<GID>166</GID>
<name>IN_1</name></connection>
<intersection>42 5</intersection>
<intersection>48 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>48,-111,48,-107.5</points>
<connection>
<GID>163</GID>
<name>N_in0</name></connection>
<intersection>-111 1</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>42,-111,42,-107.5</points>
<connection>
<GID>156</GID>
<name>nQ</name></connection>
<intersection>-111 1</intersection></vsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31,-110,31,-109</points>
<intersection>-110 2</intersection>
<intersection>-109 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31,-109,36,-109</points>
<intersection>31 0</intersection>
<intersection>36 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>29.5,-110,31,-110</points>
<connection>
<GID>166</GID>
<name>OUT</name></connection>
<intersection>31 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>36,-109,36,-107.5</points>
<connection>
<GID>156</GID>
<name>K</name></connection>
<intersection>-109 1</intersection></vsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-14,-136.5,-12.5,-136.5</points>
<connection>
<GID>169</GID>
<name>clock</name></connection>
<connection>
<GID>172</GID>
<name>CLK</name></connection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-3.5,-134.5,-3.5,-132.5</points>
<intersection>-134.5 2</intersection>
<intersection>-132.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-3.5,-132.5,-0.5,-132.5</points>
<connection>
<GID>173</GID>
<name>N_in0</name></connection>
<intersection>-3.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-6.5,-134.5,-3.5,-134.5</points>
<connection>
<GID>169</GID>
<name>Q</name></connection>
<intersection>-3.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-26,-134.5,-26,-134</points>
<connection>
<GID>170</GID>
<name>OUT_0</name></connection>
<intersection>-134.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-26,-134.5,-12.5,-134.5</points>
<connection>
<GID>169</GID>
<name>J</name></connection>
<intersection>-26 0</intersection>
<intersection>-25 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>-25,-139.5,-25,-134.5</points>
<intersection>-139.5 3</intersection>
<intersection>-134.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>-25,-139.5,-12.5,-139.5</points>
<intersection>-25 2</intersection>
<intersection>-12.5 4</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-12.5,-139.5,-12.5,-138.5</points>
<connection>
<GID>169</GID>
<name>K</name></connection>
<intersection>-139.5 3</intersection></vsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-132,54.5,-131</points>
<intersection>-132 2</intersection>
<intersection>-131 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,-131,62,-131</points>
<connection>
<GID>180</GID>
<name>IN_0</name></connection>
<intersection>54.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>47,-132,54.5,-132</points>
<connection>
<GID>178</GID>
<name>OUT</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>46.5,-142,62,-142</points>
<connection>
<GID>181</GID>
<name>IN_1</name></connection>
<connection>
<GID>179</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>68,-141,76.5,-141</points>
<connection>
<GID>184</GID>
<name>N_in0</name></connection>
<connection>
<GID>181</GID>
<name>OUT</name></connection>
<intersection>69 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>69,-141,69,-135.5</points>
<intersection>-141 1</intersection>
<intersection>-135.5 4</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>62,-135.5,69,-135.5</points>
<intersection>62 5</intersection>
<intersection>69 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>62,-135.5,62,-133</points>
<connection>
<GID>180</GID>
<name>IN_1</name></connection>
<intersection>-135.5 4</intersection></vsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>68,-132,76,-132</points>
<connection>
<GID>183</GID>
<name>N_in0</name></connection>
<connection>
<GID>180</GID>
<name>OUT</name></connection>
<intersection>68.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>68.5,-138,68.5,-132</points>
<intersection>-138 4</intersection>
<intersection>-132 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>62,-138,68.5,-138</points>
<intersection>62 5</intersection>
<intersection>68.5 3</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>62,-140,62,-138</points>
<connection>
<GID>181</GID>
<name>IN_0</name></connection>
<intersection>-138 4</intersection></vsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>40.5,-141,40.5,-133</points>
<connection>
<GID>179</GID>
<name>IN_0</name></connection>
<intersection>-137 2</intersection>
<intersection>-133 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>40.5,-133,41,-133</points>
<connection>
<GID>178</GID>
<name>IN_1</name></connection>
<intersection>40.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>38,-137,40.5,-137</points>
<connection>
<GID>185</GID>
<name>CLK</name></connection>
<intersection>40.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-131,28.5,-128</points>
<connection>
<GID>182</GID>
<name>OUT_0</name></connection>
<connection>
<GID>186</GID>
<name>IN_0</name></connection>
<intersection>-131 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28.5,-131,41,-131</points>
<connection>
<GID>178</GID>
<name>IN_0</name></connection>
<intersection>28.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>92</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>28.5,-143,28.5,-133.5</points>
<connection>
<GID>186</GID>
<name>OUT_0</name></connection>
<intersection>-143 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28.5,-143,40.5,-143</points>
<connection>
<GID>179</GID>
<name>IN_1</name></connection>
<intersection>28.5 0</intersection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,33.5808,338.954,-133.958</PageViewport></page 1>
<page 2>
<PageViewport>0,33.5808,338.954,-133.958</PageViewport></page 2>
<page 3>
<PageViewport>0,33.5808,338.954,-133.958</PageViewport></page 3>
<page 4>
<PageViewport>0,33.5808,338.954,-133.958</PageViewport></page 4>
<page 5>
<PageViewport>0,33.5808,338.954,-133.958</PageViewport></page 5>
<page 6>
<PageViewport>0,33.5808,338.954,-133.958</PageViewport></page 6>
<page 7>
<PageViewport>0,33.5808,338.954,-133.958</PageViewport></page 7>
<page 8>
<PageViewport>0,33.5808,338.954,-133.958</PageViewport></page 8>
<page 9>
<PageViewport>0,33.5808,338.954,-133.958</PageViewport></page 9></circuit>
<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>13.725,-81.2,123.075,-136.475</PageViewport>
<gate>
<ID>2</ID>
<type>AA_MUX_2x1</type>
<position>33.5,-20.5</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>3 </output>
<input>
<ID>SEL_0</ID>4 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>25,-19.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_TOGGLE</type>
<position>25,-21.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>8</ID>
<type>GA_LED</type>
<position>41,-20.5</position>
<input>
<ID>N_in0</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>33.5,-13</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_LABEL</type>
<position>22,-21.5</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>AA_LABEL</type>
<position>22,-19.5</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>AA_LABEL</type>
<position>33.5,-11</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>AE_MUX_4x1</type>
<position>35.5,-42</position>
<input>
<ID>IN_0</ID>9 </input>
<input>
<ID>IN_1</ID>8 </input>
<input>
<ID>IN_2</ID>7 </input>
<input>
<ID>IN_3</ID>6 </input>
<output>
<ID>OUT</ID>12 </output>
<input>
<ID>SEL_0</ID>11 </input>
<input>
<ID>SEL_1</ID>10 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_TOGGLE</type>
<position>25.5,-39</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>24</ID>
<type>AA_TOGGLE</type>
<position>25.5,-41</position>
<output>
<ID>OUT_0</ID>7 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_TOGGLE</type>
<position>25.5,-43</position>
<output>
<ID>OUT_0</ID>8 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_TOGGLE</type>
<position>25.5,-45</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_TOGGLE</type>
<position>35,-32.5</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_TOGGLE</type>
<position>37,-32.5</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>34</ID>
<type>GA_LED</type>
<position>45,-42</position>
<input>
<ID>N_in0</ID>12 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>AA_LABEL</type>
<position>22,-39</position>
<gparam>LABEL_TEXT D3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>AA_LABEL</type>
<position>22,-41</position>
<gparam>LABEL_TEXT D2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>40</ID>
<type>AA_LABEL</type>
<position>22,-43</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>AA_LABEL</type>
<position>22,-45</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>44</ID>
<type>AA_LABEL</type>
<position>37.5,-29.5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>46</ID>
<type>AA_LABEL</type>
<position>34.5,-29.5</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>48</ID>
<type>AA_LABEL</type>
<position>46.5,-20</position>
<gparam>LABEL_TEXT OUTPUT</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>49</ID>
<type>AA_LABEL</type>
<position>50.5,-41.5</position>
<gparam>LABEL_TEXT OUTPUT</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>51</ID>
<type>AI_MUX_8x1</type>
<position>36,-67</position>
<input>
<ID>IN_0</ID>20 </input>
<input>
<ID>IN_1</ID>19 </input>
<input>
<ID>IN_2</ID>18 </input>
<input>
<ID>IN_3</ID>17 </input>
<input>
<ID>IN_4</ID>16 </input>
<input>
<ID>IN_5</ID>15 </input>
<input>
<ID>IN_6</ID>14 </input>
<input>
<ID>IN_7</ID>13 </input>
<output>
<ID>OUT</ID>24 </output>
<input>
<ID>SEL_0</ID>23 </input>
<input>
<ID>SEL_1</ID>22 </input>
<input>
<ID>SEL_2</ID>21 </input>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 8</lparam></gate>
<gate>
<ID>53</ID>
<type>AA_TOGGLE</type>
<position>24.5,-60.5</position>
<output>
<ID>OUT_0</ID>13 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>55</ID>
<type>AA_TOGGLE</type>
<position>24.5,-62.5</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>57</ID>
<type>AA_TOGGLE</type>
<position>24.5,-64.5</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>59</ID>
<type>AA_TOGGLE</type>
<position>24.5,-66.5</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>61</ID>
<type>AA_TOGGLE</type>
<position>24.5,-68.5</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>63</ID>
<type>AA_TOGGLE</type>
<position>24.5,-70.5</position>
<output>
<ID>OUT_0</ID>18 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>65</ID>
<type>AA_TOGGLE</type>
<position>24.5,-72.5</position>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>67</ID>
<type>AA_TOGGLE</type>
<position>24.5,-74.5</position>
<output>
<ID>OUT_0</ID>20 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>69</ID>
<type>AA_TOGGLE</type>
<position>33.5,-55</position>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>71</ID>
<type>AA_TOGGLE</type>
<position>36,-55</position>
<output>
<ID>OUT_0</ID>22 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>73</ID>
<type>AA_TOGGLE</type>
<position>38.5,-55</position>
<output>
<ID>OUT_0</ID>23 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>75</ID>
<type>GA_LED</type>
<position>45,-67</position>
<input>
<ID>N_in0</ID>24 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>78</ID>
<type>AA_LABEL</type>
<position>21.5,-68.5</position>
<gparam>LABEL_TEXT D3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>79</ID>
<type>AA_LABEL</type>
<position>21.5,-70.5</position>
<gparam>LABEL_TEXT D2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>80</ID>
<type>AA_LABEL</type>
<position>21.5,-72.5</position>
<gparam>LABEL_TEXT D1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>81</ID>
<type>AA_LABEL</type>
<position>21.5,-74.5</position>
<gparam>LABEL_TEXT D0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>83</ID>
<type>AA_LABEL</type>
<position>21.5,-66.5</position>
<gparam>LABEL_TEXT D4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>85</ID>
<type>AA_LABEL</type>
<position>21.5,-64.5</position>
<gparam>LABEL_TEXT D5</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>87</ID>
<type>AA_LABEL</type>
<position>21.5,-62.5</position>
<gparam>LABEL_TEXT D6</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>89</ID>
<type>AA_LABEL</type>
<position>21.5,-60</position>
<gparam>LABEL_TEXT D7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>90</ID>
<type>AA_LABEL</type>
<position>39,-52.5</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>91</ID>
<type>AA_LABEL</type>
<position>36,-52.5</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>93</ID>
<type>AA_LABEL</type>
<position>33,-52.5</position>
<gparam>LABEL_TEXT S2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>94</ID>
<type>AA_LABEL</type>
<position>50.5,-66.5</position>
<gparam>LABEL_TEXT OUTPUT</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>108</ID>
<type>AA_TOGGLE</type>
<position>29,-88.5</position>
<output>
<ID>OUT_0</ID>41 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>110</ID>
<type>AA_TOGGLE</type>
<position>38.5,-88.5</position>
<output>
<ID>OUT_0</ID>40 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>112</ID>
<type>AA_TOGGLE</type>
<position>46.5,-88.5</position>
<output>
<ID>OUT_0</ID>39 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>114</ID>
<type>AA_TOGGLE</type>
<position>54.5,-88.5</position>
<output>
<ID>OUT_0</ID>31 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>118</ID>
<type>AA_AND4</type>
<position>68.5,-98</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>34 </input>
<input>
<ID>IN_2</ID>37 </input>
<input>
<ID>IN_3</ID>38 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>120</ID>
<type>AA_AND4</type>
<position>68.5,-108</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>39 </input>
<input>
<ID>IN_2</ID>37 </input>
<input>
<ID>IN_3</ID>38 </input>
<output>
<ID>OUT</ID>43 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>122</ID>
<type>AA_AND4</type>
<position>68.5,-118.5</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>38 </input>
<input>
<ID>IN_2</ID>40 </input>
<input>
<ID>IN_3</ID>34 </input>
<output>
<ID>OUT</ID>44 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>124</ID>
<type>AA_AND4</type>
<position>68.5,-129</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>38 </input>
<input>
<ID>IN_2</ID>40 </input>
<input>
<ID>IN_3</ID>39 </input>
<output>
<ID>OUT</ID>45 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>126</ID>
<type>AA_LABEL</type>
<position>54.5,-85</position>
<gparam>LABEL_TEXT Din</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>128</ID>
<type>AA_LABEL</type>
<position>46.5,-85</position>
<gparam>LABEL_TEXT S0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>130</ID>
<type>AA_LABEL</type>
<position>38,-85</position>
<gparam>LABEL_TEXT S1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>132</ID>
<type>AA_LABEL</type>
<position>29,-85</position>
<gparam>LABEL_TEXT S2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>134</ID>
<type>AE_SMALL_INVERTER</type>
<position>33,-94</position>
<input>
<ID>IN_0</ID>41 </input>
<output>
<ID>OUT_0</ID>38 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>136</ID>
<type>AE_SMALL_INVERTER</type>
<position>42.5,-94</position>
<input>
<ID>IN_0</ID>40 </input>
<output>
<ID>OUT_0</ID>37 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>138</ID>
<type>AE_SMALL_INVERTER</type>
<position>50.5,-94</position>
<input>
<ID>IN_0</ID>39 </input>
<output>
<ID>OUT_0</ID>34 </output>
<gparam>angle 270</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>140</ID>
<type>AA_AND4</type>
<position>68.5,-139.5</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>41 </input>
<input>
<ID>IN_2</ID>37 </input>
<input>
<ID>IN_3</ID>34 </input>
<output>
<ID>OUT</ID>46 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>142</ID>
<type>AA_AND4</type>
<position>68.5,-150</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>41 </input>
<input>
<ID>IN_2</ID>37 </input>
<input>
<ID>IN_3</ID>39 </input>
<output>
<ID>OUT</ID>47 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>144</ID>
<type>AA_AND4</type>
<position>68.5,-161</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>41 </input>
<input>
<ID>IN_2</ID>40 </input>
<input>
<ID>IN_3</ID>34 </input>
<output>
<ID>OUT</ID>48 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>146</ID>
<type>AA_AND4</type>
<position>68.5,-171.5</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>41 </input>
<input>
<ID>IN_2</ID>40 </input>
<input>
<ID>IN_3</ID>39 </input>
<output>
<ID>OUT</ID>49 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>148</ID>
<type>GA_LED</type>
<position>79,-98</position>
<input>
<ID>N_in0</ID>42 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>150</ID>
<type>GA_LED</type>
<position>79,-108</position>
<input>
<ID>N_in0</ID>43 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>152</ID>
<type>GA_LED</type>
<position>79,-118.5</position>
<input>
<ID>N_in0</ID>44 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>154</ID>
<type>GA_LED</type>
<position>79,-129</position>
<input>
<ID>N_in0</ID>45 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>155</ID>
<type>GA_LED</type>
<position>79,-139.5</position>
<input>
<ID>N_in0</ID>46 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>156</ID>
<type>GA_LED</type>
<position>79,-150</position>
<input>
<ID>N_in0</ID>47 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>157</ID>
<type>GA_LED</type>
<position>79,-161</position>
<input>
<ID>N_in0</ID>48 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>158</ID>
<type>GA_LED</type>
<position>79,-171.5</position>
<input>
<ID>N_in0</ID>49 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>160</ID>
<type>AA_LABEL</type>
<position>83.5,-97.5</position>
<gparam>LABEL_TEXT O0</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>162</ID>
<type>AA_LABEL</type>
<position>84,-108</position>
<gparam>LABEL_TEXT O1</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>164</ID>
<type>AA_LABEL</type>
<position>84,-118.5</position>
<gparam>LABEL_TEXT O2</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>166</ID>
<type>AA_LABEL</type>
<position>84,-128.5</position>
<gparam>LABEL_TEXT O3</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>168</ID>
<type>AA_LABEL</type>
<position>84,-139</position>
<gparam>LABEL_TEXT O4</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>170</ID>
<type>AA_LABEL</type>
<position>84,-149.5</position>
<gparam>LABEL_TEXT O5</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>172</ID>
<type>AA_LABEL</type>
<position>84,-160.5</position>
<gparam>LABEL_TEXT O6</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>174</ID>
<type>AA_LABEL</type>
<position>83.5,-171.5</position>
<gparam>LABEL_TEXT O7</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27,-19.5,31.5,-19.5</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27,-21.5,31.5,-21.5</points>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<connection>
<GID>6</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>35.5,-20.5,40,-20.5</points>
<connection>
<GID>8</GID>
<name>N_in0</name></connection>
<connection>
<GID>2</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-18,33.5,-15</points>
<connection>
<GID>2</GID>
<name>SEL_0</name></connection>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27.5,-39,32.5,-39</points>
<connection>
<GID>20</GID>
<name>IN_3</name></connection>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27.5,-41,32.5,-41</points>
<connection>
<GID>20</GID>
<name>IN_2</name></connection>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27.5,-43,32.5,-43</points>
<connection>
<GID>20</GID>
<name>IN_1</name></connection>
<connection>
<GID>26</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>27.5,-45,32.5,-45</points>
<connection>
<GID>20</GID>
<name>IN_0</name></connection>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35.5,-37,35.5,-35.5</points>
<connection>
<GID>20</GID>
<name>SEL_1</name></connection>
<intersection>-35.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>35,-35.5,35,-34.5</points>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection>
<intersection>-35.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>35,-35.5,35.5,-35.5</points>
<intersection>35 1</intersection>
<intersection>35.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36.5,-37,36.5,-35.5</points>
<connection>
<GID>20</GID>
<name>SEL_0</name></connection>
<intersection>-35.5 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>37,-35.5,37,-34.5</points>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection>
<intersection>-35.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>36.5,-35.5,37,-35.5</points>
<intersection>36.5 0</intersection>
<intersection>37 1</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38.5,-42,44,-42</points>
<connection>
<GID>20</GID>
<name>OUT</name></connection>
<connection>
<GID>34</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-63.5,30,-60.5</points>
<intersection>-63.5 1</intersection>
<intersection>-60.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-63.5,33,-63.5</points>
<connection>
<GID>51</GID>
<name>IN_7</name></connection>
<intersection>30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26.5,-60.5,30,-60.5</points>
<connection>
<GID>53</GID>
<name>OUT_0</name></connection>
<intersection>30 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-64.5,30,-62.5</points>
<intersection>-64.5 1</intersection>
<intersection>-62.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-64.5,33,-64.5</points>
<connection>
<GID>51</GID>
<name>IN_6</name></connection>
<intersection>30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26.5,-62.5,30,-62.5</points>
<connection>
<GID>55</GID>
<name>OUT_0</name></connection>
<intersection>30 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-65.5,30,-64.5</points>
<intersection>-65.5 1</intersection>
<intersection>-64.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-65.5,33,-65.5</points>
<connection>
<GID>51</GID>
<name>IN_5</name></connection>
<intersection>30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26.5,-64.5,30,-64.5</points>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection>
<intersection>30 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>26.5,-66.5,33,-66.5</points>
<connection>
<GID>51</GID>
<name>IN_4</name></connection>
<connection>
<GID>59</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-68.5,30,-67.5</points>
<intersection>-68.5 2</intersection>
<intersection>-67.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-67.5,33,-67.5</points>
<connection>
<GID>51</GID>
<name>IN_3</name></connection>
<intersection>30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26.5,-68.5,30,-68.5</points>
<connection>
<GID>61</GID>
<name>OUT_0</name></connection>
<intersection>30 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-70.5,30,-68.5</points>
<intersection>-70.5 2</intersection>
<intersection>-68.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-68.5,33,-68.5</points>
<connection>
<GID>51</GID>
<name>IN_2</name></connection>
<intersection>30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26.5,-70.5,30,-70.5</points>
<connection>
<GID>63</GID>
<name>OUT_0</name></connection>
<intersection>30 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-72.5,30,-69.5</points>
<intersection>-72.5 2</intersection>
<intersection>-69.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-69.5,33,-69.5</points>
<connection>
<GID>51</GID>
<name>IN_1</name></connection>
<intersection>30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26.5,-72.5,30,-72.5</points>
<connection>
<GID>65</GID>
<name>OUT_0</name></connection>
<intersection>30 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>30,-74.5,30,-70.5</points>
<intersection>-74.5 2</intersection>
<intersection>-70.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-70.5,33,-70.5</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>30 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>26.5,-74.5,30,-74.5</points>
<connection>
<GID>67</GID>
<name>OUT_0</name></connection>
<intersection>30 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-61.5,35,-59</points>
<connection>
<GID>51</GID>
<name>SEL_2</name></connection>
<intersection>-59 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>33.5,-59,33.5,-57</points>
<connection>
<GID>69</GID>
<name>OUT_0</name></connection>
<intersection>-59 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>33.5,-59,35,-59</points>
<intersection>33.5 1</intersection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>36,-61.5,36,-57</points>
<connection>
<GID>51</GID>
<name>SEL_1</name></connection>
<connection>
<GID>71</GID>
<name>OUT_0</name></connection></vsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>37,-61.5,37,-59</points>
<connection>
<GID>51</GID>
<name>SEL_0</name></connection>
<intersection>-59 2</intersection></vsegment>
<vsegment>
<ID>1</ID>
<points>38.5,-59,38.5,-57</points>
<connection>
<GID>73</GID>
<name>OUT_0</name></connection>
<intersection>-59 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>37,-59,38.5,-59</points>
<intersection>37 0</intersection>
<intersection>38.5 1</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>39,-67,44,-67</points>
<connection>
<GID>51</GID>
<name>OUT</name></connection>
<connection>
<GID>75</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54.5,-168.5,54.5,-90.5</points>
<connection>
<GID>114</GID>
<name>OUT_0</name></connection>
<intersection>-168.5 15</intersection>
<intersection>-158 13</intersection>
<intersection>-147 11</intersection>
<intersection>-136.5 9</intersection>
<intersection>-126 7</intersection>
<intersection>-115.5 5</intersection>
<intersection>-105 3</intersection>
<intersection>-95 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54.5,-95,65.5,-95</points>
<connection>
<GID>118</GID>
<name>IN_0</name></connection>
<intersection>54.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>54.5,-105,65.5,-105</points>
<connection>
<GID>120</GID>
<name>IN_0</name></connection>
<intersection>54.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>54.5,-115.5,65.5,-115.5</points>
<connection>
<GID>122</GID>
<name>IN_0</name></connection>
<intersection>54.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>54.5,-126,65.5,-126</points>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<intersection>54.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>54.5,-136.5,65.5,-136.5</points>
<connection>
<GID>140</GID>
<name>IN_0</name></connection>
<intersection>54.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>54.5,-147,65.5,-147</points>
<connection>
<GID>142</GID>
<name>IN_0</name></connection>
<intersection>54.5 0</intersection></hsegment>
<hsegment>
<ID>13</ID>
<points>54.5,-158,65.5,-158</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<intersection>54.5 0</intersection></hsegment>
<hsegment>
<ID>15</ID>
<points>54.5,-168.5,65.5,-168.5</points>
<connection>
<GID>146</GID>
<name>IN_0</name></connection>
<intersection>54.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-164,50.5,-96</points>
<connection>
<GID>138</GID>
<name>OUT_0</name></connection>
<intersection>-164 7</intersection>
<intersection>-142.5 5</intersection>
<intersection>-121.5 3</intersection>
<intersection>-97 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50.5,-97,65.5,-97</points>
<connection>
<GID>118</GID>
<name>IN_1</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>50.5,-121.5,65.5,-121.5</points>
<connection>
<GID>122</GID>
<name>IN_3</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>50.5,-142.5,65.5,-142.5</points>
<connection>
<GID>140</GID>
<name>IN_3</name></connection>
<intersection>50.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>50.5,-164,65.5,-164</points>
<connection>
<GID>144</GID>
<name>IN_3</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>42.5,-151,42.5,-96</points>
<connection>
<GID>136</GID>
<name>OUT_0</name></connection>
<intersection>-151 9</intersection>
<intersection>-140.5 7</intersection>
<intersection>-109 3</intersection>
<intersection>-99 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42.5,-99,65.5,-99</points>
<connection>
<GID>118</GID>
<name>IN_2</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>42.5,-109,65.5,-109</points>
<connection>
<GID>120</GID>
<name>IN_2</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>42.5,-140.5,65.5,-140.5</points>
<connection>
<GID>140</GID>
<name>IN_2</name></connection>
<intersection>42.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>42.5,-151,65.5,-151</points>
<connection>
<GID>142</GID>
<name>IN_2</name></connection>
<intersection>42.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-128,33,-96</points>
<connection>
<GID>134</GID>
<name>OUT_0</name></connection>
<intersection>-128 7</intersection>
<intersection>-117.5 5</intersection>
<intersection>-111 3</intersection>
<intersection>-101 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33,-101,65.5,-101</points>
<connection>
<GID>118</GID>
<name>IN_3</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>33,-111,65.5,-111</points>
<connection>
<GID>120</GID>
<name>IN_3</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>33,-117.5,65.5,-117.5</points>
<connection>
<GID>122</GID>
<name>IN_1</name></connection>
<intersection>33 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>33,-128,65.5,-128</points>
<connection>
<GID>124</GID>
<name>IN_1</name></connection>
<intersection>33 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>46.5,-174.5,46.5,-90.5</points>
<connection>
<GID>112</GID>
<name>OUT_0</name></connection>
<intersection>-174.5 7</intersection>
<intersection>-153 5</intersection>
<intersection>-132 3</intersection>
<intersection>-107 1</intersection>
<intersection>-92 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>46.5,-107,65.5,-107</points>
<connection>
<GID>120</GID>
<name>IN_1</name></connection>
<intersection>46.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>46.5,-132,65.5,-132</points>
<connection>
<GID>124</GID>
<name>IN_3</name></connection>
<intersection>46.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>46.5,-153,65.5,-153</points>
<connection>
<GID>142</GID>
<name>IN_3</name></connection>
<intersection>46.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>46.5,-174.5,65.5,-174.5</points>
<connection>
<GID>146</GID>
<name>IN_3</name></connection>
<intersection>46.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>46.5,-92,50.5,-92</points>
<connection>
<GID>138</GID>
<name>IN_0</name></connection>
<intersection>46.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-172.5,38.5,-90.5</points>
<connection>
<GID>110</GID>
<name>OUT_0</name></connection>
<intersection>-172.5 7</intersection>
<intersection>-162 5</intersection>
<intersection>-130 3</intersection>
<intersection>-119.5 1</intersection>
<intersection>-92 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38.5,-119.5,65.5,-119.5</points>
<connection>
<GID>122</GID>
<name>IN_2</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>38.5,-130,65.5,-130</points>
<connection>
<GID>124</GID>
<name>IN_2</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>38.5,-162,65.5,-162</points>
<connection>
<GID>144</GID>
<name>IN_2</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>38.5,-172.5,65.5,-172.5</points>
<connection>
<GID>146</GID>
<name>IN_2</name></connection>
<intersection>38.5 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>38.5,-92,42.5,-92</points>
<connection>
<GID>136</GID>
<name>IN_0</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>29,-170.5,29,-90.5</points>
<connection>
<GID>108</GID>
<name>OUT_0</name></connection>
<intersection>-170.5 7</intersection>
<intersection>-160 5</intersection>
<intersection>-149 3</intersection>
<intersection>-138.5 1</intersection>
<intersection>-92 8</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>29,-138.5,65.5,-138.5</points>
<connection>
<GID>140</GID>
<name>IN_1</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>29,-149,65.5,-149</points>
<connection>
<GID>142</GID>
<name>IN_1</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>29,-160,65.5,-160</points>
<connection>
<GID>144</GID>
<name>IN_1</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>29,-170.5,65.5,-170.5</points>
<connection>
<GID>146</GID>
<name>IN_1</name></connection>
<intersection>29 0</intersection></hsegment>
<hsegment>
<ID>8</ID>
<points>29,-92,33,-92</points>
<connection>
<GID>134</GID>
<name>IN_0</name></connection>
<intersection>29 0</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71.5,-98,78,-98</points>
<connection>
<GID>118</GID>
<name>OUT</name></connection>
<connection>
<GID>148</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71.5,-108,78,-108</points>
<connection>
<GID>150</GID>
<name>N_in0</name></connection>
<connection>
<GID>120</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71.5,-118.5,78,-118.5</points>
<connection>
<GID>152</GID>
<name>N_in0</name></connection>
<connection>
<GID>122</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71.5,-129,78,-129</points>
<connection>
<GID>154</GID>
<name>N_in0</name></connection>
<connection>
<GID>124</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71.5,-139.5,78,-139.5</points>
<connection>
<GID>155</GID>
<name>N_in0</name></connection>
<connection>
<GID>140</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71.5,-150,78,-150</points>
<connection>
<GID>142</GID>
<name>OUT</name></connection>
<connection>
<GID>156</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71.5,-161,78,-161</points>
<connection>
<GID>144</GID>
<name>OUT</name></connection>
<connection>
<GID>157</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>71.5,-171.5,78,-171.5</points>
<connection>
<GID>146</GID>
<name>OUT</name></connection>
<connection>
<GID>158</GID>
<name>N_in0</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 1>
<page 2>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 2>
<page 3>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 3>
<page 4>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 4>
<page 5>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 5>
<page 6>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 6>
<page 7>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 7>
<page 8>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 8>
<page 9>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 9></circuit>
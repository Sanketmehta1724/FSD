<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-535.743,-329.918,-248.394,-475.17</PageViewport>
<gate>
<ID>194</ID>
<type>AA_LABEL</type>
<position>-461,-118.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>195</ID>
<type>AA_LABEL</type>
<position>-442,-118.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>199</ID>
<type>BA_NAND2</type>
<position>-435.5,-127</position>
<input>
<ID>IN_0</ID>85 </input>
<input>
<ID>IN_1</ID>85 </input>
<output>
<ID>OUT</ID>83 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>201</ID>
<type>BA_NAND2</type>
<position>-420.5,-140</position>
<input>
<ID>IN_0</ID>89 </input>
<input>
<ID>IN_1</ID>83 </input>
<output>
<ID>OUT</ID>86 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>203</ID>
<type>BA_NAND2</type>
<position>-420,-149</position>
<input>
<ID>IN_0</ID>84 </input>
<input>
<ID>IN_1</ID>85 </input>
<output>
<ID>OUT</ID>87 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>205</ID>
<type>BA_NAND2</type>
<position>-403,-144.5</position>
<input>
<ID>IN_0</ID>86 </input>
<input>
<ID>IN_1</ID>87 </input>
<output>
<ID>OUT</ID>88 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>12</ID>
<type>BA_NAND2</type>
<position>-400,191.5</position>
<input>
<ID>IN_0</ID>1 </input>
<output>
<ID>OUT</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>207</ID>
<type>GA_LED</type>
<position>-391,-144.5</position>
<input>
<ID>N_in0</ID>88 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>AA_TOGGLE</type>
<position>-409.5,191.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>209</ID>
<type>BA_NAND2</type>
<position>-421.5,-160.5</position>
<input>
<ID>IN_0</ID>89 </input>
<input>
<ID>IN_1</ID>85 </input>
<output>
<ID>OUT</ID>90 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>16</ID>
<type>GA_LED</type>
<position>-388.5,191.5</position>
<input>
<ID>N_in0</ID>2 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>211</ID>
<type>BA_NAND2</type>
<position>-407,-160.5</position>
<input>
<ID>IN_0</ID>90 </input>
<input>
<ID>IN_1</ID>90 </input>
<output>
<ID>OUT</ID>91 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_LABEL</type>
<position>-397,198.5</position>
<gparam>LABEL_TEXT Nand As A Not Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>212</ID>
<type>GA_LED</type>
<position>-394.5,-160.5</position>
<input>
<ID>N_in0</ID>91 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>214</ID>
<type>AA_LABEL</type>
<position>-390,-140</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>216</ID>
<type>AA_LABEL</type>
<position>-392.5,-155.5</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>217</ID>
<type>AA_LABEL</type>
<position>-433.5,-178</position>
<gparam>LABEL_TEXT __________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>218</ID>
<type>AA_LABEL</type>
<position>-428.5,-185.5</position>
<gparam>LABEL_TEXT Half-subtractor</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>219</ID>
<type>AA_AND2</type>
<position>-426,-226</position>
<input>
<ID>IN_0</ID>101 </input>
<input>
<ID>IN_1</ID>94 </input>
<output>
<ID>OUT</ID>96 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>26</ID>
<type>BA_NAND2</type>
<position>-400,179.5</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>5 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>220</ID>
<type>AA_AND2</type>
<position>-426,-231.5</position>
<input>
<ID>IN_0</ID>95 </input>
<input>
<ID>IN_1</ID>93 </input>
<output>
<ID>OUT</ID>97 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>221</ID>
<type>AA_AND2</type>
<position>-425.5,-238.5</position>
<input>
<ID>IN_0</ID>95 </input>
<input>
<ID>IN_1</ID>93 </input>
<output>
<ID>OUT</ID>99 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>222</ID>
<type>AA_TOGGLE</type>
<position>-457,-206.5</position>
<output>
<ID>OUT_0</ID>101 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>223</ID>
<type>AA_TOGGLE</type>
<position>-444,-206.5</position>
<output>
<ID>OUT_0</ID>93 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_TOGGLE</type>
<position>-410,181</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>224</ID>
<type>AE_SMALL_INVERTER</type>
<position>-453,-210.5</position>
<input>
<ID>IN_0</ID>101 </input>
<output>
<ID>OUT_0</ID>95 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>225</ID>
<type>AE_SMALL_INVERTER</type>
<position>-440.5,-210</position>
<input>
<ID>IN_0</ID>93 </input>
<output>
<ID>OUT_0</ID>94 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_TOGGLE</type>
<position>-410,178.5</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>226</ID>
<type>AE_OR2</type>
<position>-414,-228</position>
<input>
<ID>IN_0</ID>96 </input>
<input>
<ID>IN_1</ID>97 </input>
<output>
<ID>OUT</ID>98 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>227</ID>
<type>GA_LED</type>
<position>-404,-227.5</position>
<input>
<ID>N_in0</ID>98 </input>
<input>
<ID>N_in1</ID>100 </input>
<input>
<ID>N_in2</ID>100 </input>
<input>
<ID>N_in3</ID>100 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>228</ID>
<type>GA_LED</type>
<position>-416,-238.5</position>
<input>
<ID>N_in0</ID>99 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>AA_LABEL</type>
<position>-398,186</position>
<gparam>LABEL_TEXT Nand As And Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>229</ID>
<type>AA_LABEL</type>
<position>-444,-200</position>
<gparam>LABEL_TEXT AOI Implementation</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>BA_NAND2</type>
<position>-390,179.5</position>
<input>
<ID>IN_0</ID>8 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>230</ID>
<type>AI_XOR2</type>
<position>-344.5,-211</position>
<input>
<ID>IN_0</ID>106 </input>
<input>
<ID>IN_1</ID>103 </input>
<output>
<ID>OUT</ID>104 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>37</ID>
<type>GA_LED</type>
<position>-382.5,179.5</position>
<input>
<ID>N_in0</ID>9 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>231</ID>
<type>AA_AND2</type>
<position>-344,-220.5</position>
<input>
<ID>IN_0</ID>107 </input>
<input>
<ID>IN_1</ID>103 </input>
<output>
<ID>OUT</ID>105 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>38</ID>
<type>BA_NAND2</type>
<position>-400.5,163.5</position>
<input>
<ID>IN_0</ID>10 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>232</ID>
<type>AA_TOGGLE</type>
<position>-359.5,-214.5</position>
<output>
<ID>OUT_0</ID>106 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>39</ID>
<type>BA_NAND2</type>
<position>-400,156</position>
<input>
<ID>IN_0</ID>11 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>233</ID>
<type>AA_TOGGLE</type>
<position>-359,-216.5</position>
<output>
<ID>OUT_0</ID>103 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>40</ID>
<type>AA_TOGGLE</type>
<position>-408.5,163.5</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>234</ID>
<type>GA_LED</type>
<position>-335.5,-211</position>
<input>
<ID>N_in0</ID>104 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>41</ID>
<type>AA_TOGGLE</type>
<position>-408.5,156.5</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>235</ID>
<type>GA_LED</type>
<position>-335.5,-220</position>
<input>
<ID>N_in0</ID>105 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>236</ID>
<type>AA_LABEL</type>
<position>-404,-223</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>237</ID>
<type>AA_LABEL</type>
<position>-416.5,-234.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>44</ID>
<type>BA_NAND2</type>
<position>-387.5,160</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>13 </input>
<output>
<ID>OUT</ID>20 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>45</ID>
<type>GA_LED</type>
<position>-377.5,160</position>
<input>
<ID>N_in0</ID>20 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>46</ID>
<type>AA_LABEL</type>
<position>-397.5,170.5</position>
<gparam>LABEL_TEXT Nand As Or Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>240</ID>
<type>AE_SMALL_INVERTER</type>
<position>-348.5,-215.5</position>
<input>
<ID>IN_0</ID>106 </input>
<output>
<ID>OUT_0</ID>107 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>47</ID>
<type>BA_NAND2</type>
<position>-401,139.5</position>
<input>
<ID>IN_0</ID>15 </input>
<output>
<ID>OUT</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>241</ID>
<type>AA_LABEL</type>
<position>-472.5,-274.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>48</ID>
<type>BA_NAND2</type>
<position>-400.5,132</position>
<input>
<ID>IN_0</ID>16 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>242</ID>
<type>AA_LABEL</type>
<position>-453.5,-274.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>49</ID>
<type>AA_TOGGLE</type>
<position>-409.5,139.5</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>243</ID>
<type>BA_NAND2</type>
<position>-447,-283</position>
<input>
<ID>IN_0</ID>110 </input>
<input>
<ID>IN_1</ID>110 </input>
<output>
<ID>OUT</ID>108 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>50</ID>
<type>AA_TOGGLE</type>
<position>-410.5,131</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>244</ID>
<type>BA_NAND2</type>
<position>-432,-296</position>
<input>
<ID>IN_0</ID>117 </input>
<input>
<ID>IN_1</ID>108 </input>
<output>
<ID>OUT</ID>111 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>51</ID>
<type>BA_NAND2</type>
<position>-388,136</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>18 </input>
<output>
<ID>OUT</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>245</ID>
<type>BA_NAND2</type>
<position>-431.5,-305</position>
<input>
<ID>IN_0</ID>109 </input>
<input>
<ID>IN_1</ID>110 </input>
<output>
<ID>OUT</ID>112 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>246</ID>
<type>BA_NAND2</type>
<position>-414.5,-300.5</position>
<input>
<ID>IN_0</ID>111 </input>
<input>
<ID>IN_1</ID>112 </input>
<output>
<ID>OUT</ID>113 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>53</ID>
<type>AA_LABEL</type>
<position>-398,146.5</position>
<gparam>LABEL_TEXT Nand As Nor Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>247</ID>
<type>GA_LED</type>
<position>-402.5,-300.5</position>
<input>
<ID>N_in0</ID>113 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>54</ID>
<type>BA_NAND2</type>
<position>-376,136.5</position>
<input>
<ID>IN_0</ID>21 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>248</ID>
<type>BA_NAND2</type>
<position>-433,-316.5</position>
<input>
<ID>IN_0</ID>109 </input>
<input>
<ID>IN_1</ID>110 </input>
<output>
<ID>OUT</ID>115 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>249</ID>
<type>BA_NAND2</type>
<position>-418.5,-316.5</position>
<input>
<ID>IN_0</ID>115 </input>
<input>
<ID>IN_1</ID>115 </input>
<output>
<ID>OUT</ID>116 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>56</ID>
<type>GA_LED</type>
<position>-366.5,136.5</position>
<input>
<ID>N_in0</ID>22 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>250</ID>
<type>GA_LED</type>
<position>-406,-316.5</position>
<input>
<ID>N_in0</ID>116 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>251</ID>
<type>AA_LABEL</type>
<position>-401.5,-296</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>58</ID>
<type>BA_NAND2</type>
<position>-400,112.5</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>25 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>252</ID>
<type>AA_LABEL</type>
<position>-404,-311.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>253</ID>
<type>AA_LABEL</type>
<position>-458,-269.5</position>
<gparam>LABEL_TEXT Nand Implementation</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>BA_NAND2</type>
<position>-388,120.5</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>25 </input>
<output>
<ID>OUT</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>254</ID>
<type>AA_TOGGLE</type>
<position>-472.5,-277.5</position>
<output>
<ID>OUT_0</ID>117 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>255</ID>
<type>AA_TOGGLE</type>
<position>-453.5,-277.5</position>
<output>
<ID>OUT_0</ID>110 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>62</ID>
<type>BA_NAND2</type>
<position>-389,106.5</position>
<input>
<ID>IN_0</ID>25 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>256</ID>
<type>BA_NAND2</type>
<position>-466.5,-283</position>
<input>
<ID>IN_0</ID>117 </input>
<input>
<ID>IN_1</ID>117 </input>
<output>
<ID>OUT</ID>109 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>257</ID>
<type>AA_LABEL</type>
<position>-441.5,-346</position>
<gparam>LABEL_TEXT __________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>64</ID>
<type>BA_NAND2</type>
<position>-375,114</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>28 </input>
<output>
<ID>OUT</ID>29 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>258</ID>
<type>AA_LABEL</type>
<position>-421,-354.5</position>
<gparam>LABEL_TEXT Full-Adder</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>259</ID>
<type>AA_LABEL</type>
<position>-464.5,-362.5</position>
<gparam>LABEL_TEXT Nand Implementation</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>66</ID>
<type>AA_TOGGLE</type>
<position>-410.5,120</position>
<output>
<ID>OUT_0</ID>23 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>261</ID>
<type>AA_TOGGLE</type>
<position>-473.5,-370.5</position>
<output>
<ID>OUT_0</ID>126 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>68</ID>
<type>AA_TOGGLE</type>
<position>-410.5,105</position>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>263</ID>
<type>AA_TOGGLE</type>
<position>-450,-370.5</position>
<output>
<ID>OUT_0</ID>124 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>70</ID>
<type>GA_LED</type>
<position>-361,114</position>
<input>
<ID>N_in0</ID>29 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>71</ID>
<type>AA_LABEL</type>
<position>-396.5,126.5</position>
<gparam>LABEL_TEXT Nand As Xor Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>265</ID>
<type>AA_TOGGLE</type>
<position>-429.5,-370.5</position>
<output>
<ID>OUT_0</ID>122 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>72</ID>
<type>BA_NAND2</type>
<position>-400,79</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>73</ID>
<type>BA_NAND2</type>
<position>-388,87</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>31 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>267</ID>
<type>BA_NAND2</type>
<position>-463.5,-383.5</position>
<input>
<ID>IN_0</ID>126 </input>
<input>
<ID>IN_1</ID>126 </input>
<output>
<ID>OUT</ID>120 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>74</ID>
<type>BA_NAND2</type>
<position>-389,73</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>34 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>75</ID>
<type>BA_NAND2</type>
<position>-375,78.5</position>
<input>
<ID>IN_0</ID>33 </input>
<input>
<ID>IN_1</ID>34 </input>
<output>
<ID>OUT</ID>39 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>269</ID>
<type>BA_NAND2</type>
<position>-439.5,-383.5</position>
<input>
<ID>IN_0</ID>124 </input>
<input>
<ID>IN_1</ID>124 </input>
<output>
<ID>OUT</ID>121 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>76</ID>
<type>AA_TOGGLE</type>
<position>-410.5,86.5</position>
<output>
<ID>OUT_0</ID>30 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>77</ID>
<type>AA_TOGGLE</type>
<position>-410,71</position>
<output>
<ID>OUT_0</ID>32 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>271</ID>
<type>BA_NAND2</type>
<position>-418,-383</position>
<input>
<ID>IN_0</ID>122 </input>
<input>
<ID>IN_1</ID>122 </input>
<output>
<ID>OUT</ID>125 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>79</ID>
<type>AA_LABEL</type>
<position>-396.5,93</position>
<gparam>LABEL_TEXT Nand As Xnor Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>80</ID>
<type>BA_NAND2</type>
<position>-361.5,78.5</position>
<input>
<ID>IN_0</ID>39 </input>
<input>
<ID>IN_1</ID>39 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>81</ID>
<type>GA_LED</type>
<position>-350.5,78.5</position>
<input>
<ID>N_in0</ID>40 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>83</ID>
<type>AA_LABEL</type>
<position>-417,87</position>
<gparam>LABEL_TEXT input-a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>84</ID>
<type>AA_LABEL</type>
<position>-416,121</position>
<gparam>LABEL_TEXT input-a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>85</ID>
<type>AA_LABEL</type>
<position>-415,140</position>
<gparam>LABEL_TEXT input-a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>86</ID>
<type>AA_LABEL</type>
<position>-414.5,164</position>
<gparam>LABEL_TEXT input-a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>87</ID>
<type>AA_LABEL</type>
<position>-415,181.5</position>
<gparam>LABEL_TEXT input-a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>88</ID>
<type>AA_LABEL</type>
<position>-414.5,192.5</position>
<gparam>LABEL_TEXT input-a</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>90</ID>
<type>AA_LABEL</type>
<position>-415.5,179</position>
<gparam>LABEL_TEXT input-b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>91</ID>
<type>AA_LABEL</type>
<position>-414,156.5</position>
<gparam>LABEL_TEXT input-b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>92</ID>
<type>AA_LABEL</type>
<position>-415,131.5</position>
<gparam>LABEL_TEXT input-b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>93</ID>
<type>AA_LABEL</type>
<position>-415,105.5</position>
<gparam>LABEL_TEXT input-b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>94</ID>
<type>AA_LABEL</type>
<position>-416.5,71.5</position>
<gparam>LABEL_TEXT input-b</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>289</ID>
<type>BA_NAND3</type>
<position>-399,-392.5</position>
<input>
<ID>IN_0</ID>120 </input>
<input>
<ID>IN_1</ID>121 </input>
<input>
<ID>IN_2</ID>122 </input>
<output>
<ID>OUT</ID>131 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>291</ID>
<type>BA_NAND3</type>
<position>-399,-401.5</position>
<input>
<ID>IN_0</ID>120 </input>
<input>
<ID>IN_1</ID>124 </input>
<input>
<ID>IN_2</ID>125 </input>
<output>
<ID>OUT</ID>132 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>98</ID>
<type>AA_LABEL</type>
<position>-427.5,63</position>
<gparam>LABEL_TEXT __________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________________</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>99</ID>
<type>AA_LABEL</type>
<position>-393.5,56</position>
<gparam>LABEL_TEXT Nor As A Not Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>293</ID>
<type>BA_NAND3</type>
<position>-399,-410</position>
<input>
<ID>IN_0</ID>126 </input>
<input>
<ID>IN_1</ID>121 </input>
<input>
<ID>IN_2</ID>125 </input>
<output>
<ID>OUT</ID>133 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>101</ID>
<type>BE_NOR2</type>
<position>-396,47.5</position>
<input>
<ID>IN_0</ID>41 </input>
<input>
<ID>IN_1</ID>41 </input>
<output>
<ID>OUT</ID>42 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>295</ID>
<type>BA_NAND3</type>
<position>-399,-419</position>
<input>
<ID>IN_0</ID>126 </input>
<input>
<ID>IN_1</ID>124 </input>
<input>
<ID>IN_2</ID>122 </input>
<output>
<ID>OUT</ID>134 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>103</ID>
<type>AA_TOGGLE</type>
<position>-403.5,48</position>
<output>
<ID>OUT_0</ID>41 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>297</ID>
<type>BA_NAND3</type>
<position>-398.5,-448</position>
<input>
<ID>IN_0</ID>126 </input>
<input>
<ID>IN_1</ID>121 </input>
<input>
<ID>IN_2</ID>122 </input>
<output>
<ID>OUT</ID>136 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>105</ID>
<type>GA_LED</type>
<position>-386,47.5</position>
<input>
<ID>N_in0</ID>42 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>299</ID>
<type>BA_NAND3</type>
<position>-398.5,-439</position>
<input>
<ID>IN_0</ID>120 </input>
<input>
<ID>IN_1</ID>124 </input>
<input>
<ID>IN_2</ID>122 </input>
<output>
<ID>OUT</ID>135 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>106</ID>
<type>AA_LABEL</type>
<position>-393.5,21</position>
<gparam>LABEL_TEXT Nor As A Xnor Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>301</ID>
<type>BA_NAND3</type>
<position>-398.5,-457</position>
<input>
<ID>IN_0</ID>126 </input>
<input>
<ID>IN_1</ID>124 </input>
<input>
<ID>IN_2</ID>125 </input>
<output>
<ID>OUT</ID>137 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>108</ID>
<type>BE_NOR2</type>
<position>-399.5,10</position>
<input>
<ID>IN_0</ID>43 </input>
<input>
<ID>IN_1</ID>44 </input>
<output>
<ID>OUT</ID>45 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>303</ID>
<type>BA_NAND3</type>
<position>-398.5,-466.5</position>
<input>
<ID>IN_0</ID>126 </input>
<input>
<ID>IN_1</ID>124 </input>
<input>
<ID>IN_2</ID>122 </input>
<output>
<ID>OUT</ID>138 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 3</lparam></gate>
<gate>
<ID>110</ID>
<type>BE_NOR2</type>
<position>-390,15.5</position>
<input>
<ID>IN_0</ID>43 </input>
<input>
<ID>IN_1</ID>45 </input>
<output>
<ID>OUT</ID>46 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>112</ID>
<type>BE_NOR2</type>
<position>-389.5,5</position>
<input>
<ID>IN_0</ID>45 </input>
<input>
<ID>IN_1</ID>44 </input>
<output>
<ID>OUT</ID>47 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>307</ID>
<type>BA_NAND4</type>
<position>-363.5,-452.5</position>
<input>
<ID>IN_0</ID>135 </input>
<input>
<ID>IN_1</ID>136 </input>
<input>
<ID>IN_2</ID>137 </input>
<input>
<ID>IN_3</ID>138 </input>
<output>
<ID>OUT</ID>141 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>114</ID>
<type>BE_NOR2</type>
<position>-378.5,10.5</position>
<input>
<ID>IN_0</ID>46 </input>
<input>
<ID>IN_1</ID>47 </input>
<output>
<ID>OUT</ID>48 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>309</ID>
<type>BA_NAND4</type>
<position>-361,-404.5</position>
<input>
<ID>IN_0</ID>131 </input>
<input>
<ID>IN_1</ID>132 </input>
<input>
<ID>IN_2</ID>133 </input>
<input>
<ID>IN_3</ID>134 </input>
<output>
<ID>OUT</ID>139 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 4</lparam></gate>
<gate>
<ID>116</ID>
<type>AA_TOGGLE</type>
<position>-411,16</position>
<output>
<ID>OUT_0</ID>43 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>311</ID>
<type>GA_LED</type>
<position>-339.5,-404.5</position>
<input>
<ID>N_in0</ID>139 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>118</ID>
<type>AA_TOGGLE</type>
<position>-411,5.5</position>
<output>
<ID>OUT_0</ID>44 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>120</ID>
<type>GA_LED</type>
<position>-368.5,10.5</position>
<input>
<ID>N_in0</ID>48 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>121</ID>
<type>AA_LABEL</type>
<position>-395.5,42.5</position>
<gparam>LABEL_TEXT Nor As A Xor Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>122</ID>
<type>BE_NOR2</type>
<position>-401.5,31.5</position>
<input>
<ID>IN_0</ID>49 </input>
<input>
<ID>IN_1</ID>50 </input>
<output>
<ID>OUT</ID>51 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>123</ID>
<type>BE_NOR2</type>
<position>-392,37</position>
<input>
<ID>IN_0</ID>49 </input>
<input>
<ID>IN_1</ID>51 </input>
<output>
<ID>OUT</ID>52 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>317</ID>
<type>GA_LED</type>
<position>-349,-452.5</position>
<input>
<ID>N_in0</ID>141 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>124</ID>
<type>BE_NOR2</type>
<position>-391.5,26.5</position>
<input>
<ID>IN_0</ID>51 </input>
<input>
<ID>IN_1</ID>50 </input>
<output>
<ID>OUT</ID>53 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>318</ID>
<type>AA_LABEL</type>
<position>-339.5,-399.5</position>
<gparam>LABEL_TEXT S</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>125</ID>
<type>BE_NOR2</type>
<position>-380.5,32</position>
<input>
<ID>IN_0</ID>52 </input>
<input>
<ID>IN_1</ID>53 </input>
<output>
<ID>OUT</ID>55 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>319</ID>
<type>AA_LABEL</type>
<position>-349.5,-448</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>126</ID>
<type>AA_TOGGLE</type>
<position>-413,37.5</position>
<output>
<ID>OUT_0</ID>49 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>320</ID>
<type>AA_LABEL</type>
<position>-450.5,-365.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>127</ID>
<type>AA_TOGGLE</type>
<position>-413,27</position>
<output>
<ID>OUT_0</ID>50 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>321</ID>
<type>AA_LABEL</type>
<position>-473.5,-366</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>128</ID>
<type>GA_LED</type>
<position>-359.5,31.5</position>
<input>
<ID>N_in0</ID>56 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>322</ID>
<type>AA_LABEL</type>
<position>-429.5,-365</position>
<gparam>LABEL_TEXT C</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>129</ID>
<type>BE_NOR2</type>
<position>-370,31.5</position>
<input>
<ID>IN_0</ID>55 </input>
<input>
<ID>IN_1</ID>55 </input>
<output>
<ID>OUT</ID>56 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>131</ID>
<type>AA_TOGGLE</type>
<position>-409,-12</position>
<output>
<ID>OUT_0</ID>58 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>133</ID>
<type>BE_NOR2</type>
<position>-393.5,-13</position>
<input>
<ID>IN_0</ID>58 </input>
<input>
<ID>IN_1</ID>59 </input>
<output>
<ID>OUT</ID>57 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>135</ID>
<type>BE_NOR2</type>
<position>-376.5,-13</position>
<input>
<ID>IN_0</ID>57 </input>
<input>
<ID>IN_1</ID>57 </input>
<output>
<ID>OUT</ID>60 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>136</ID>
<type>AA_TOGGLE</type>
<position>-409,-14</position>
<output>
<ID>OUT_0</ID>59 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>137</ID>
<type>GA_LED</type>
<position>-367,-13</position>
<input>
<ID>N_in0</ID>60 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>138</ID>
<type>AA_LABEL</type>
<position>-393,-4.5</position>
<gparam>LABEL_TEXT Nor As A Or Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>139</ID>
<type>BE_NOR2</type>
<position>-398,-29.5</position>
<input>
<ID>IN_0</ID>61 </input>
<input>
<ID>IN_1</ID>61 </input>
<output>
<ID>OUT</ID>63 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>140</ID>
<type>BE_NOR2</type>
<position>-398,-39</position>
<input>
<ID>IN_0</ID>62 </input>
<input>
<ID>IN_1</ID>62 </input>
<output>
<ID>OUT</ID>64 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>141</ID>
<type>BE_NOR2</type>
<position>-385.5,-33.5</position>
<input>
<ID>IN_0</ID>63 </input>
<input>
<ID>IN_1</ID>64 </input>
<output>
<ID>OUT</ID>65 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>142</ID>
<type>AA_TOGGLE</type>
<position>-407.5,-29.5</position>
<output>
<ID>OUT_0</ID>61 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>143</ID>
<type>AA_TOGGLE</type>
<position>-407,-38.5</position>
<output>
<ID>OUT_0</ID>62 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>144</ID>
<type>GA_LED</type>
<position>-375,-33</position>
<input>
<ID>N_in0</ID>65 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>145</ID>
<type>AA_LABEL</type>
<position>-391.5,-22.5</position>
<gparam>LABEL_TEXT Nor As A AND Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>147</ID>
<type>AA_LABEL</type>
<position>-380,-51.5</position>
<gparam>LABEL_TEXT Half-Adder</gparam>
<gparam>TEXT_HEIGHT 4</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>149</ID>
<type>AA_AND2</type>
<position>-409,-86.5</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>70 </input>
<output>
<ID>OUT</ID>72 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>151</ID>
<type>AA_AND2</type>
<position>-409,-92</position>
<input>
<ID>IN_0</ID>71 </input>
<input>
<ID>IN_1</ID>69 </input>
<output>
<ID>OUT</ID>73 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>153</ID>
<type>AA_AND2</type>
<position>-408.5,-99</position>
<input>
<ID>IN_0</ID>68 </input>
<input>
<ID>IN_1</ID>69 </input>
<output>
<ID>OUT</ID>75 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>157</ID>
<type>AA_TOGGLE</type>
<position>-440,-67</position>
<output>
<ID>OUT_0</ID>68 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>159</ID>
<type>AA_TOGGLE</type>
<position>-427,-67</position>
<output>
<ID>OUT_0</ID>69 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>161</ID>
<type>AE_SMALL_INVERTER</type>
<position>-436,-71</position>
<input>
<ID>IN_0</ID>68 </input>
<output>
<ID>OUT_0</ID>71 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>163</ID>
<type>AE_SMALL_INVERTER</type>
<position>-423.5,-70.5</position>
<input>
<ID>IN_0</ID>69 </input>
<output>
<ID>OUT_0</ID>70 </output>
<gparam>angle 0.0</gparam>
<lparam>DEFAULT_DELAY 1</lparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>165</ID>
<type>AE_OR2</type>
<position>-397,-88.5</position>
<input>
<ID>IN_0</ID>72 </input>
<input>
<ID>IN_1</ID>73 </input>
<output>
<ID>OUT</ID>74 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>167</ID>
<type>GA_LED</type>
<position>-387,-88</position>
<input>
<ID>N_in0</ID>74 </input>
<input>
<ID>N_in1</ID>76 </input>
<input>
<ID>N_in2</ID>76 </input>
<input>
<ID>N_in3</ID>76 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>169</ID>
<type>GA_LED</type>
<position>-399,-99</position>
<input>
<ID>N_in0</ID>75 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>171</ID>
<type>AA_LABEL</type>
<position>-427,-60.5</position>
<gparam>LABEL_TEXT AOI Implementation</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>173</ID>
<type>AI_XOR2</type>
<position>-334,-78.5</position>
<input>
<ID>IN_0</ID>77 </input>
<input>
<ID>IN_1</ID>79 </input>
<output>
<ID>OUT</ID>80 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>175</ID>
<type>AA_AND2</type>
<position>-333.5,-88</position>
<input>
<ID>IN_0</ID>77 </input>
<input>
<ID>IN_1</ID>79 </input>
<output>
<ID>OUT</ID>81 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>177</ID>
<type>AA_TOGGLE</type>
<position>-349,-82</position>
<output>
<ID>OUT_0</ID>77 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>179</ID>
<type>AA_TOGGLE</type>
<position>-349,-84</position>
<output>
<ID>OUT_0</ID>79 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>181</ID>
<type>GA_LED</type>
<position>-325,-78.5</position>
<input>
<ID>N_in0</ID>80 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>183</ID>
<type>GA_LED</type>
<position>-325,-87.5</position>
<input>
<ID>N_in0</ID>81 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>184</ID>
<type>AA_LABEL</type>
<position>-446.5,-113.5</position>
<gparam>LABEL_TEXT Nand Implementation</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>186</ID>
<type>AA_TOGGLE</type>
<position>-461,-121.5</position>
<output>
<ID>OUT_0</ID>89 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>188</ID>
<type>AA_TOGGLE</type>
<position>-442,-121.5</position>
<output>
<ID>OUT_0</ID>85 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>192</ID>
<type>BA_NAND2</type>
<position>-455,-127</position>
<input>
<ID>IN_0</ID>89 </input>
<input>
<ID>IN_1</ID>89 </input>
<output>
<ID>OUT</ID>84 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-407.5,190.5,-403,190.5</points>
<intersection>-407.5 3</intersection>
<intersection>-403 4</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-407.5,190.5,-407.5,191.5</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>190.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>-403,190.5,-403,192.5</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>190.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-397,191.5,-389.5,191.5</points>
<connection>
<GID>12</GID>
<name>OUT</name></connection>
<connection>
<GID>16</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-408,178.5,-403,178.5</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<connection>
<GID>32</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-405.5,180.5,-405.5,181</points>
<intersection>180.5 1</intersection>
<intersection>181 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-405.5,180.5,-403,180.5</points>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>-405.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-408,181,-405.5,181</points>
<connection>
<GID>30</GID>
<name>OUT_0</name></connection>
<intersection>-405.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-393,178.5,-393,180.5</points>
<connection>
<GID>36</GID>
<name>IN_0</name></connection>
<intersection>178.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-397,178.5,-393,178.5</points>
<intersection>-397 3</intersection>
<intersection>-393 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-397,178.5,-397,179.5</points>
<connection>
<GID>26</GID>
<name>OUT</name></connection>
<intersection>178.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-387,179.5,-383.5,179.5</points>
<connection>
<GID>37</GID>
<name>N_in0</name></connection>
<connection>
<GID>36</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-403.5,162.5,-403.5,164.5</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>162.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-406.5,162.5,-403.5,162.5</points>
<intersection>-406.5 3</intersection>
<intersection>-403.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-406.5,162.5,-406.5,163.5</points>
<connection>
<GID>40</GID>
<name>OUT_0</name></connection>
<intersection>162.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-402.5,155,-402.5,157</points>
<intersection>155 2</intersection>
<intersection>157 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-403,157,-402.5,157</points>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>-402.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-406.5,155,-402.5,155</points>
<intersection>-406.5 3</intersection>
<intersection>-402.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-406.5,155,-406.5,156.5</points>
<connection>
<GID>41</GID>
<name>OUT_0</name></connection>
<intersection>155 2</intersection></vsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-394,161,-394,163.5</points>
<intersection>161 1</intersection>
<intersection>163.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-394,161,-390.5,161</points>
<connection>
<GID>44</GID>
<name>IN_0</name></connection>
<intersection>-394 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-397.5,163.5,-394,163.5</points>
<connection>
<GID>38</GID>
<name>OUT</name></connection>
<intersection>-394 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-393.5,156,-393.5,159</points>
<intersection>156 2</intersection>
<intersection>159 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-393.5,159,-390.5,159</points>
<connection>
<GID>44</GID>
<name>IN_1</name></connection>
<intersection>-393.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-397,156,-393.5,156</points>
<connection>
<GID>39</GID>
<name>OUT</name></connection>
<intersection>-393.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-404,139.5,-404,140.5</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<intersection>139.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-407.5,139.5,-404,139.5</points>
<connection>
<GID>49</GID>
<name>OUT_0</name></connection>
<intersection>-404 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-403,131,-403,133</points>
<intersection>131 2</intersection>
<intersection>133 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-403.5,133,-403,133</points>
<connection>
<GID>48</GID>
<name>IN_0</name></connection>
<intersection>-403 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-408.5,131,-403,131</points>
<connection>
<GID>50</GID>
<name>OUT_0</name></connection>
<intersection>-403 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-394.5,137,-394.5,139.5</points>
<intersection>137 1</intersection>
<intersection>139.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-394.5,137,-391,137</points>
<connection>
<GID>51</GID>
<name>IN_0</name></connection>
<intersection>-394.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-398,139.5,-394.5,139.5</points>
<connection>
<GID>47</GID>
<name>OUT</name></connection>
<intersection>-394.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-394,132,-394,135</points>
<intersection>132 2</intersection>
<intersection>135 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-394,135,-391,135</points>
<connection>
<GID>51</GID>
<name>IN_1</name></connection>
<intersection>-394 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-397.5,132,-394,132</points>
<connection>
<GID>48</GID>
<name>OUT</name></connection>
<intersection>-394 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-384.5,160,-378.5,160</points>
<connection>
<GID>45</GID>
<name>N_in0</name></connection>
<connection>
<GID>44</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-382,135.5,-382,136</points>
<intersection>135.5 1</intersection>
<intersection>136 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-382,135.5,-379,135.5</points>
<intersection>-382 0</intersection>
<intersection>-379 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-385,136,-382,136</points>
<connection>
<GID>51</GID>
<name>OUT</name></connection>
<intersection>-382 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-379,135.5,-379,137.5</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>135.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-373,136.5,-367.5,136.5</points>
<connection>
<GID>56</GID>
<name>N_in0</name></connection>
<connection>
<GID>54</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-403.5,113.5,-403.5,120.5</points>
<intersection>113.5 1</intersection>
<intersection>120.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-403.5,113.5,-403,113.5</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>-403.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-408.5,120.5,-391,120.5</points>
<intersection>-408.5 3</intersection>
<intersection>-403.5 0</intersection>
<intersection>-391 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-408.5,120,-408.5,120.5</points>
<connection>
<GID>66</GID>
<name>OUT_0</name></connection>
<intersection>120.5 2</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-391,120.5,-391,121.5</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>120.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-394.5,107.5,-394.5,119.5</points>
<intersection>107.5 3</intersection>
<intersection>112.5 1</intersection>
<intersection>119.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-397,112.5,-394.5,112.5</points>
<connection>
<GID>58</GID>
<name>OUT</name></connection>
<intersection>-394.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-394.5,119.5,-391,119.5</points>
<connection>
<GID>60</GID>
<name>IN_1</name></connection>
<intersection>-394.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-394.5,107.5,-392,107.5</points>
<connection>
<GID>62</GID>
<name>IN_0</name></connection>
<intersection>-394.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-408.5,105,-392,105</points>
<connection>
<GID>68</GID>
<name>OUT_0</name></connection>
<intersection>-403 4</intersection>
<intersection>-392 11</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-403,105,-403,111.5</points>
<connection>
<GID>58</GID>
<name>IN_1</name></connection>
<intersection>105 1</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>-392,105,-392,105.5</points>
<connection>
<GID>62</GID>
<name>IN_1</name></connection>
<intersection>105 1</intersection></vsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-380.5,115,-380.5,120.5</points>
<intersection>115 1</intersection>
<intersection>120.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-380.5,115,-378,115</points>
<connection>
<GID>64</GID>
<name>IN_0</name></connection>
<intersection>-380.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-385,120.5,-380.5,120.5</points>
<connection>
<GID>60</GID>
<name>OUT</name></connection>
<intersection>-380.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-380.5,106.5,-380.5,113</points>
<intersection>106.5 1</intersection>
<intersection>113 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-386,106.5,-380.5,106.5</points>
<connection>
<GID>62</GID>
<name>OUT</name></connection>
<intersection>-380.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-380.5,113,-378,113</points>
<connection>
<GID>64</GID>
<name>IN_1</name></connection>
<intersection>-380.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<hsegment>
<ID>2</ID>
<points>-372,114,-362,114</points>
<connection>
<GID>64</GID>
<name>OUT</name></connection>
<connection>
<GID>70</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-403.5,80,-403.5,87</points>
<intersection>80 1</intersection>
<intersection>87 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-403.5,80,-403,80</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<intersection>-403.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-408.5,87,-391,87</points>
<intersection>-408.5 3</intersection>
<intersection>-403.5 0</intersection>
<intersection>-391 5</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-408.5,86.5,-408.5,87</points>
<connection>
<GID>76</GID>
<name>OUT_0</name></connection>
<intersection>87 2</intersection></vsegment>
<vsegment>
<ID>5</ID>
<points>-391,87,-391,88</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>87 2</intersection></vsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-394.5,74,-394.5,86</points>
<intersection>74 3</intersection>
<intersection>79 1</intersection>
<intersection>86 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-397,79,-394.5,79</points>
<connection>
<GID>72</GID>
<name>OUT</name></connection>
<intersection>-394.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-394.5,86,-391,86</points>
<connection>
<GID>73</GID>
<name>IN_1</name></connection>
<intersection>-394.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-394.5,74,-392,74</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>-394.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-408,71,-392,71</points>
<connection>
<GID>77</GID>
<name>OUT_0</name></connection>
<intersection>-403 4</intersection>
<intersection>-392 11</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>-403,71,-403,78</points>
<connection>
<GID>72</GID>
<name>IN_1</name></connection>
<intersection>71 1</intersection></vsegment>
<vsegment>
<ID>11</ID>
<points>-392,71,-392,72</points>
<connection>
<GID>74</GID>
<name>IN_1</name></connection>
<intersection>71 1</intersection></vsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-380.5,79.5,-380.5,87</points>
<intersection>79.5 1</intersection>
<intersection>87 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-380.5,79.5,-378,79.5</points>
<connection>
<GID>75</GID>
<name>IN_0</name></connection>
<intersection>-380.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-385,87,-380.5,87</points>
<connection>
<GID>73</GID>
<name>OUT</name></connection>
<intersection>-380.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-380.5,73,-380.5,77.5</points>
<intersection>73 1</intersection>
<intersection>77.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-386,73,-380.5,73</points>
<connection>
<GID>74</GID>
<name>OUT</name></connection>
<intersection>-380.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-380.5,77.5,-378,77.5</points>
<connection>
<GID>75</GID>
<name>IN_1</name></connection>
<intersection>-380.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-368,78,-368,78.5</points>
<intersection>78 1</intersection>
<intersection>78.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-368,78,-364.5,78</points>
<intersection>-368 0</intersection>
<intersection>-364.5 3</intersection>
<intersection>-364.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-372,78.5,-368,78.5</points>
<connection>
<GID>75</GID>
<name>OUT</name></connection>
<intersection>-368 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-364.5,77.5,-364.5,79.5</points>
<connection>
<GID>80</GID>
<name>IN_0</name></connection>
<connection>
<GID>80</GID>
<name>IN_1</name></connection>
<intersection>78 1</intersection></vsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-358.5,78.5,-351.5,78.5</points>
<connection>
<GID>81</GID>
<name>N_in0</name></connection>
<connection>
<GID>80</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-399.5,48,-399.5,48.5</points>
<intersection>48 2</intersection>
<intersection>48.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-399.5,48.5,-398,48.5</points>
<connection>
<GID>101</GID>
<name>IN_0</name></connection>
<intersection>-399.5 0</intersection>
<intersection>-398 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-401.5,48,-399.5,48</points>
<connection>
<GID>103</GID>
<name>OUT_0</name></connection>
<intersection>-399.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-398,46.5,-398,48.5</points>
<intersection>46.5 4</intersection>
<intersection>48.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-399,46.5,-398,46.5</points>
<connection>
<GID>101</GID>
<name>IN_1</name></connection>
<intersection>-398 3</intersection></hsegment></shape></wire>
<wire>
<ID>42</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-393,47.5,-387,47.5</points>
<connection>
<GID>101</GID>
<name>OUT</name></connection>
<connection>
<GID>105</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>43</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-401,16,-401,16.5</points>
<intersection>16 2</intersection>
<intersection>16.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-401,16.5,-393,16.5</points>
<connection>
<GID>110</GID>
<name>IN_0</name></connection>
<intersection>-401 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-409,16,-401,16</points>
<connection>
<GID>116</GID>
<name>OUT_0</name></connection>
<intersection>-402.5 3</intersection>
<intersection>-401 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-402.5,11,-402.5,16</points>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<intersection>16 2</intersection></vsegment></shape></wire>
<wire>
<ID>44</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-400.5,4,-400.5,5.5</points>
<intersection>4 1</intersection>
<intersection>5.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-400.5,4,-392.5,4</points>
<connection>
<GID>112</GID>
<name>IN_1</name></connection>
<intersection>-400.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-409,5.5,-400.5,5.5</points>
<connection>
<GID>118</GID>
<name>OUT_0</name></connection>
<intersection>-402.5 3</intersection>
<intersection>-400.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-402.5,5.5,-402.5,9</points>
<connection>
<GID>108</GID>
<name>IN_1</name></connection>
<intersection>5.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>45</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-394.5,6,-394.5,14.5</points>
<intersection>6 3</intersection>
<intersection>10 1</intersection>
<intersection>14.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-396.5,10,-394.5,10</points>
<connection>
<GID>108</GID>
<name>OUT</name></connection>
<intersection>-394.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-394.5,14.5,-393,14.5</points>
<connection>
<GID>110</GID>
<name>IN_1</name></connection>
<intersection>-394.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-394.5,6,-392.5,6</points>
<connection>
<GID>112</GID>
<name>IN_0</name></connection>
<intersection>-394.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>46</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-384,11.5,-384,15.5</points>
<intersection>11.5 1</intersection>
<intersection>15.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-384,11.5,-381.5,11.5</points>
<connection>
<GID>114</GID>
<name>IN_0</name></connection>
<intersection>-384 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-387,15.5,-384,15.5</points>
<connection>
<GID>110</GID>
<name>OUT</name></connection>
<intersection>-384 0</intersection></hsegment></shape></wire>
<wire>
<ID>47</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-384,5,-384,9.5</points>
<intersection>5 1</intersection>
<intersection>9.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-386.5,5,-384,5</points>
<connection>
<GID>112</GID>
<name>OUT</name></connection>
<intersection>-384 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-384,9.5,-381.5,9.5</points>
<connection>
<GID>114</GID>
<name>IN_1</name></connection>
<intersection>-384 0</intersection></hsegment></shape></wire>
<wire>
<ID>48</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-375.5,10.5,-369.5,10.5</points>
<connection>
<GID>120</GID>
<name>N_in0</name></connection>
<connection>
<GID>114</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>49</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-403,37.5,-403,38</points>
<intersection>37.5 2</intersection>
<intersection>38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-403,38,-395,38</points>
<connection>
<GID>123</GID>
<name>IN_0</name></connection>
<intersection>-403 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-411,37.5,-403,37.5</points>
<connection>
<GID>126</GID>
<name>OUT_0</name></connection>
<intersection>-404.5 3</intersection>
<intersection>-403 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-404.5,32.5,-404.5,37.5</points>
<connection>
<GID>122</GID>
<name>IN_0</name></connection>
<intersection>37.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>50</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-402.5,25.5,-402.5,27</points>
<intersection>25.5 1</intersection>
<intersection>27 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-402.5,25.5,-394.5,25.5</points>
<connection>
<GID>124</GID>
<name>IN_1</name></connection>
<intersection>-402.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-411,27,-402.5,27</points>
<connection>
<GID>127</GID>
<name>OUT_0</name></connection>
<intersection>-404.5 3</intersection>
<intersection>-402.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-404.5,27,-404.5,30.5</points>
<connection>
<GID>122</GID>
<name>IN_1</name></connection>
<intersection>27 2</intersection></vsegment></shape></wire>
<wire>
<ID>51</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-396.5,27.5,-396.5,36</points>
<intersection>27.5 3</intersection>
<intersection>31.5 1</intersection>
<intersection>36 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-398.5,31.5,-396.5,31.5</points>
<connection>
<GID>122</GID>
<name>OUT</name></connection>
<intersection>-396.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-396.5,36,-395,36</points>
<connection>
<GID>123</GID>
<name>IN_1</name></connection>
<intersection>-396.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-396.5,27.5,-394.5,27.5</points>
<connection>
<GID>124</GID>
<name>IN_0</name></connection>
<intersection>-396.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>52</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-386,33,-386,37</points>
<intersection>33 1</intersection>
<intersection>37 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-386,33,-383.5,33</points>
<connection>
<GID>125</GID>
<name>IN_0</name></connection>
<intersection>-386 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-389,37,-386,37</points>
<connection>
<GID>123</GID>
<name>OUT</name></connection>
<intersection>-386 0</intersection></hsegment></shape></wire>
<wire>
<ID>53</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-386,26.5,-386,31</points>
<intersection>26.5 1</intersection>
<intersection>31 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-388.5,26.5,-386,26.5</points>
<connection>
<GID>124</GID>
<name>OUT</name></connection>
<intersection>-386 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-386,31,-383.5,31</points>
<connection>
<GID>125</GID>
<name>IN_1</name></connection>
<intersection>-386 0</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-377.5,32.5,-373,32.5</points>
<connection>
<GID>129</GID>
<name>IN_0</name></connection>
<intersection>-377.5 6</intersection>
<intersection>-374 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-374,30.5,-374,32.5</points>
<intersection>30.5 4</intersection>
<intersection>32.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-374,30.5,-373,30.5</points>
<connection>
<GID>129</GID>
<name>IN_1</name></connection>
<intersection>-374 3</intersection></hsegment>
<vsegment>
<ID>6</ID>
<points>-377.5,32,-377.5,32.5</points>
<connection>
<GID>125</GID>
<name>OUT</name></connection>
<intersection>32.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-367,31.5,-360.5,31.5</points>
<connection>
<GID>129</GID>
<name>OUT</name></connection>
<connection>
<GID>128</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-385,-13,-385,-12</points>
<intersection>-13 1</intersection>
<intersection>-12 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-390.5,-13,-385,-13</points>
<connection>
<GID>133</GID>
<name>OUT</name></connection>
<intersection>-385 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-385,-12,-379.5,-12</points>
<connection>
<GID>135</GID>
<name>IN_0</name></connection>
<intersection>-385 0</intersection>
<intersection>-380.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-380.5,-14,-380.5,-12</points>
<intersection>-14 4</intersection>
<intersection>-12 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>-380.5,-14,-379.5,-14</points>
<connection>
<GID>135</GID>
<name>IN_1</name></connection>
<intersection>-380.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-407,-12,-396.5,-12</points>
<connection>
<GID>131</GID>
<name>OUT_0</name></connection>
<connection>
<GID>133</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-407,-14,-396.5,-14</points>
<connection>
<GID>133</GID>
<name>IN_1</name></connection>
<connection>
<GID>136</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-373.5,-13,-368,-13</points>
<connection>
<GID>135</GID>
<name>OUT</name></connection>
<connection>
<GID>137</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-403,-29.5,-403,-28.5</points>
<intersection>-29.5 2</intersection>
<intersection>-28.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-403,-28.5,-401,-28.5</points>
<connection>
<GID>139</GID>
<name>IN_0</name></connection>
<intersection>-403 0</intersection>
<intersection>-401 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-405.5,-29.5,-403,-29.5</points>
<connection>
<GID>142</GID>
<name>OUT_0</name></connection>
<intersection>-403 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-401,-30.5,-401,-28.5</points>
<connection>
<GID>139</GID>
<name>IN_1</name></connection>
<intersection>-28.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-403,-38.5,-403,-38</points>
<intersection>-38.5 6</intersection>
<intersection>-38 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-403,-38,-401,-38</points>
<connection>
<GID>140</GID>
<name>IN_0</name></connection>
<intersection>-403 0</intersection>
<intersection>-401 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-401,-40,-401,-38</points>
<connection>
<GID>140</GID>
<name>IN_1</name></connection>
<intersection>-38 2</intersection></vsegment>
<hsegment>
<ID>6</ID>
<points>-405,-38.5,-403,-38.5</points>
<connection>
<GID>143</GID>
<name>OUT_0</name></connection>
<intersection>-403 0</intersection></hsegment></shape></wire>
<wire>
<ID>63</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-391.5,-32.5,-391.5,-29.5</points>
<intersection>-32.5 2</intersection>
<intersection>-29.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-395,-29.5,-391.5,-29.5</points>
<connection>
<GID>139</GID>
<name>OUT</name></connection>
<intersection>-391.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-391.5,-32.5,-388.5,-32.5</points>
<connection>
<GID>141</GID>
<name>IN_0</name></connection>
<intersection>-391.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>64</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-391.5,-39,-391.5,-34.5</points>
<intersection>-39 1</intersection>
<intersection>-34.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-395,-39,-391.5,-39</points>
<connection>
<GID>140</GID>
<name>OUT</name></connection>
<intersection>-391.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-391.5,-34.5,-388.5,-34.5</points>
<connection>
<GID>141</GID>
<name>IN_1</name></connection>
<intersection>-391.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>65</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-379,-33.5,-379,-33</points>
<intersection>-33.5 2</intersection>
<intersection>-33 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-379,-33,-376,-33</points>
<connection>
<GID>144</GID>
<name>N_in0</name></connection>
<intersection>-379 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-382.5,-33.5,-379,-33.5</points>
<connection>
<GID>141</GID>
<name>OUT</name></connection>
<intersection>-379 0</intersection></hsegment></shape></wire>
<wire>
<ID>68</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-440,-98,-440,-69</points>
<connection>
<GID>157</GID>
<name>OUT_0</name></connection>
<intersection>-98 4</intersection>
<intersection>-85.5 1</intersection>
<intersection>-71 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-440,-85.5,-412,-85.5</points>
<connection>
<GID>149</GID>
<name>IN_0</name></connection>
<intersection>-440 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-440,-71,-438,-71</points>
<connection>
<GID>161</GID>
<name>IN_0</name></connection>
<intersection>-440 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-440,-98,-411.5,-98</points>
<connection>
<GID>153</GID>
<name>IN_0</name></connection>
<intersection>-440 0</intersection></hsegment></shape></wire>
<wire>
<ID>69</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-427,-100,-427,-69</points>
<connection>
<GID>159</GID>
<name>OUT_0</name></connection>
<intersection>-100 4</intersection>
<intersection>-93 1</intersection>
<intersection>-70.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-427,-93,-412,-93</points>
<connection>
<GID>151</GID>
<name>IN_1</name></connection>
<intersection>-427 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-427,-70.5,-425.5,-70.5</points>
<connection>
<GID>163</GID>
<name>IN_0</name></connection>
<intersection>-427 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-427,-100,-411.5,-100</points>
<connection>
<GID>153</GID>
<name>IN_1</name></connection>
<intersection>-427 0</intersection></hsegment></shape></wire>
<wire>
<ID>70</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-416.5,-87.5,-416.5,-70.5</points>
<intersection>-87.5 1</intersection>
<intersection>-70.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-416.5,-87.5,-412,-87.5</points>
<connection>
<GID>149</GID>
<name>IN_1</name></connection>
<intersection>-416.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-421.5,-70.5,-416.5,-70.5</points>
<connection>
<GID>163</GID>
<name>OUT_0</name></connection>
<intersection>-416.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>71</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-423,-91,-423,-71</points>
<intersection>-91 1</intersection>
<intersection>-71 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-423,-91,-412,-91</points>
<connection>
<GID>151</GID>
<name>IN_0</name></connection>
<intersection>-423 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-434,-71,-423,-71</points>
<connection>
<GID>161</GID>
<name>OUT_0</name></connection>
<intersection>-423 0</intersection></hsegment></shape></wire>
<wire>
<ID>72</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-402.5,-87.5,-402.5,-86.5</points>
<intersection>-87.5 1</intersection>
<intersection>-86.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-402.5,-87.5,-400,-87.5</points>
<connection>
<GID>165</GID>
<name>IN_0</name></connection>
<intersection>-402.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-406,-86.5,-402.5,-86.5</points>
<connection>
<GID>149</GID>
<name>OUT</name></connection>
<intersection>-402.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-403,-92,-403,-89.5</points>
<intersection>-92 2</intersection>
<intersection>-89.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-403,-89.5,-400,-89.5</points>
<connection>
<GID>165</GID>
<name>IN_1</name></connection>
<intersection>-403 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-406,-92,-403,-92</points>
<connection>
<GID>151</GID>
<name>OUT</name></connection>
<intersection>-403 0</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-391,-88.5,-391,-88</points>
<intersection>-88.5 2</intersection>
<intersection>-88 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-391,-88,-388,-88</points>
<connection>
<GID>167</GID>
<name>N_in0</name></connection>
<intersection>-391 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-394,-88.5,-391,-88.5</points>
<connection>
<GID>165</GID>
<name>OUT</name></connection>
<intersection>-391 0</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-405.5,-99,-400,-99</points>
<connection>
<GID>153</GID>
<name>OUT</name></connection>
<connection>
<GID>169</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-387,-89,-387,-87</points>
<connection>
<GID>167</GID>
<name>N_in3</name></connection>
<connection>
<GID>167</GID>
<name>N_in2</name></connection>
<intersection>-88 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-387,-88,-386,-88</points>
<connection>
<GID>167</GID>
<name>N_in1</name></connection>
<intersection>-387 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-339,-87,-339,-77.5</points>
<intersection>-87 5</intersection>
<intersection>-82 2</intersection>
<intersection>-77.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-339,-77.5,-337,-77.5</points>
<connection>
<GID>173</GID>
<name>IN_0</name></connection>
<intersection>-339 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-347,-82,-339,-82</points>
<connection>
<GID>177</GID>
<name>OUT_0</name></connection>
<intersection>-339 0</intersection></hsegment>
<hsegment>
<ID>5</ID>
<points>-339,-87,-336.5,-87</points>
<connection>
<GID>175</GID>
<name>IN_0</name></connection>
<intersection>-339 0</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-341.5,-89,-341.5,-79.5</points>
<intersection>-89 1</intersection>
<intersection>-84 2</intersection>
<intersection>-79.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-341.5,-89,-336.5,-89</points>
<connection>
<GID>175</GID>
<name>IN_1</name></connection>
<intersection>-341.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-347,-84,-341.5,-84</points>
<connection>
<GID>179</GID>
<name>OUT_0</name></connection>
<intersection>-341.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-341.5,-79.5,-337,-79.5</points>
<connection>
<GID>173</GID>
<name>IN_1</name></connection>
<intersection>-341.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-331,-78.5,-326,-78.5</points>
<connection>
<GID>181</GID>
<name>N_in0</name></connection>
<connection>
<GID>173</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-328,-88,-328,-87.5</points>
<intersection>-88 2</intersection>
<intersection>-87.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-328,-87.5,-326,-87.5</points>
<connection>
<GID>183</GID>
<name>N_in0</name></connection>
<intersection>-328 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-330.5,-88,-328,-88</points>
<connection>
<GID>175</GID>
<name>OUT</name></connection>
<intersection>-328 0</intersection></hsegment></shape></wire>
<wire>
<ID>83</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-428,-141,-428,-127</points>
<intersection>-141 1</intersection>
<intersection>-127 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-428,-141,-423.5,-141</points>
<connection>
<GID>201</GID>
<name>IN_1</name></connection>
<intersection>-428 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-432.5,-127,-428,-127</points>
<connection>
<GID>199</GID>
<name>OUT</name></connection>
<intersection>-428 0</intersection></hsegment></shape></wire>
<wire>
<ID>84</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-452.5,-148,-452.5,-127</points>
<intersection>-148 2</intersection>
<intersection>-127 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-452.5,-127,-452,-127</points>
<connection>
<GID>192</GID>
<name>OUT</name></connection>
<intersection>-452.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-452.5,-148,-423,-148</points>
<connection>
<GID>203</GID>
<name>IN_0</name></connection>
<intersection>-452.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>85</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-442,-161.5,-442,-123.5</points>
<connection>
<GID>188</GID>
<name>OUT_0</name></connection>
<intersection>-161.5 14</intersection>
<intersection>-150 8</intersection>
<intersection>-127 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-442,-127,-438.5,-127</points>
<intersection>-442 0</intersection>
<intersection>-438.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-438.5,-128,-438.5,-126</points>
<connection>
<GID>199</GID>
<name>IN_1</name></connection>
<connection>
<GID>199</GID>
<name>IN_0</name></connection>
<intersection>-127 2</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-442,-150,-423,-150</points>
<connection>
<GID>203</GID>
<name>IN_1</name></connection>
<intersection>-442 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>-442,-161.5,-424.5,-161.5</points>
<connection>
<GID>209</GID>
<name>IN_1</name></connection>
<intersection>-442 0</intersection></hsegment></shape></wire>
<wire>
<ID>86</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-411.5,-143.5,-411.5,-140</points>
<intersection>-143.5 1</intersection>
<intersection>-140 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-411.5,-143.5,-406,-143.5</points>
<connection>
<GID>205</GID>
<name>IN_0</name></connection>
<intersection>-411.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-417.5,-140,-411.5,-140</points>
<connection>
<GID>201</GID>
<name>OUT</name></connection>
<intersection>-411.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>87</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-411.5,-149,-411.5,-145.5</points>
<intersection>-149 2</intersection>
<intersection>-145.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-411.5,-145.5,-406,-145.5</points>
<connection>
<GID>205</GID>
<name>IN_1</name></connection>
<intersection>-411.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-417,-149,-411.5,-149</points>
<connection>
<GID>203</GID>
<name>OUT</name></connection>
<intersection>-411.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>88</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-400,-144.5,-392,-144.5</points>
<connection>
<GID>207</GID>
<name>N_in0</name></connection>
<intersection>-400 11</intersection></hsegment>
<vsegment>
<ID>11</ID>
<points>-400,-144.5,-400,-144.5</points>
<connection>
<GID>205</GID>
<name>OUT</name></connection>
<intersection>-144.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>89</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-461,-159.5,-461,-123.5</points>
<connection>
<GID>186</GID>
<name>OUT_0</name></connection>
<intersection>-159.5 1</intersection>
<intersection>-139 3</intersection>
<intersection>-127 4</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-461,-159.5,-424.5,-159.5</points>
<connection>
<GID>209</GID>
<name>IN_0</name></connection>
<intersection>-461 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-461,-139,-423.5,-139</points>
<connection>
<GID>201</GID>
<name>IN_0</name></connection>
<intersection>-461 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-461,-127,-458,-127</points>
<intersection>-461 0</intersection>
<intersection>-458 5</intersection></hsegment>
<vsegment>
<ID>5</ID>
<points>-458,-128,-458,-126</points>
<connection>
<GID>192</GID>
<name>IN_1</name></connection>
<connection>
<GID>192</GID>
<name>IN_0</name></connection>
<intersection>-127 4</intersection></vsegment></shape></wire>
<wire>
<ID>90</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-418.5,-160.5,-410,-160.5</points>
<connection>
<GID>209</GID>
<name>OUT</name></connection>
<intersection>-410 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-410,-161.5,-410,-159.5</points>
<connection>
<GID>211</GID>
<name>IN_1</name></connection>
<connection>
<GID>211</GID>
<name>IN_0</name></connection>
<intersection>-160.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>91</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-404,-160.5,-395.5,-160.5</points>
<connection>
<GID>212</GID>
<name>N_in0</name></connection>
<connection>
<GID>211</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>93</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-444,-239.5,-444,-208.5</points>
<connection>
<GID>223</GID>
<name>OUT_0</name></connection>
<intersection>-239.5 4</intersection>
<intersection>-232.5 1</intersection>
<intersection>-210 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-444,-232.5,-429,-232.5</points>
<connection>
<GID>220</GID>
<name>IN_1</name></connection>
<intersection>-444 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-444,-210,-442.5,-210</points>
<connection>
<GID>225</GID>
<name>IN_0</name></connection>
<intersection>-444 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-444,-239.5,-428.5,-239.5</points>
<connection>
<GID>221</GID>
<name>IN_1</name></connection>
<intersection>-444 0</intersection></hsegment></shape></wire>
<wire>
<ID>94</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-433.5,-227,-433.5,-210</points>
<intersection>-227 1</intersection>
<intersection>-210 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-433.5,-227,-429,-227</points>
<connection>
<GID>219</GID>
<name>IN_1</name></connection>
<intersection>-433.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-438.5,-210,-433.5,-210</points>
<connection>
<GID>225</GID>
<name>OUT_0</name></connection>
<intersection>-433.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>95</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-451,-237.5,-451,-210.5</points>
<connection>
<GID>224</GID>
<name>OUT_0</name></connection>
<intersection>-237.5 3</intersection>
<intersection>-230.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-451,-230.5,-429,-230.5</points>
<connection>
<GID>220</GID>
<name>IN_0</name></connection>
<intersection>-451 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-451,-237.5,-428.5,-237.5</points>
<connection>
<GID>221</GID>
<name>IN_0</name></connection>
<intersection>-451 0</intersection></hsegment></shape></wire>
<wire>
<ID>96</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-419.5,-227,-419.5,-226</points>
<intersection>-227 1</intersection>
<intersection>-226 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-419.5,-227,-417,-227</points>
<connection>
<GID>226</GID>
<name>IN_0</name></connection>
<intersection>-419.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-423,-226,-419.5,-226</points>
<connection>
<GID>219</GID>
<name>OUT</name></connection>
<intersection>-419.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>97</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-420,-231.5,-420,-229</points>
<intersection>-231.5 2</intersection>
<intersection>-229 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-420,-229,-417,-229</points>
<connection>
<GID>226</GID>
<name>IN_1</name></connection>
<intersection>-420 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-423,-231.5,-420,-231.5</points>
<connection>
<GID>220</GID>
<name>OUT</name></connection>
<intersection>-420 0</intersection></hsegment></shape></wire>
<wire>
<ID>98</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-408,-228,-408,-227.5</points>
<intersection>-228 2</intersection>
<intersection>-227.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-408,-227.5,-405,-227.5</points>
<connection>
<GID>227</GID>
<name>N_in0</name></connection>
<intersection>-408 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-411,-228,-408,-228</points>
<connection>
<GID>226</GID>
<name>OUT</name></connection>
<intersection>-408 0</intersection></hsegment></shape></wire>
<wire>
<ID>99</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-422.5,-238.5,-417,-238.5</points>
<connection>
<GID>228</GID>
<name>N_in0</name></connection>
<connection>
<GID>221</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>100</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-404,-228.5,-404,-226.5</points>
<connection>
<GID>227</GID>
<name>N_in3</name></connection>
<connection>
<GID>227</GID>
<name>N_in2</name></connection>
<intersection>-227.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-404,-227.5,-403,-227.5</points>
<connection>
<GID>227</GID>
<name>N_in1</name></connection>
<intersection>-404 0</intersection></hsegment></shape></wire>
<wire>
<ID>101</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-457,-225,-457,-208.5</points>
<connection>
<GID>222</GID>
<name>OUT_0</name></connection>
<intersection>-225 1</intersection>
<intersection>-210.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-457,-225,-429,-225</points>
<connection>
<GID>219</GID>
<name>IN_0</name></connection>
<intersection>-457 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-457,-210.5,-455,-210.5</points>
<connection>
<GID>224</GID>
<name>IN_0</name></connection>
<intersection>-457 0</intersection></hsegment></shape></wire>
<wire>
<ID>103</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-352,-221.5,-352,-212</points>
<intersection>-221.5 1</intersection>
<intersection>-216.5 2</intersection>
<intersection>-212 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-352,-221.5,-347,-221.5</points>
<connection>
<GID>231</GID>
<name>IN_1</name></connection>
<intersection>-352 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-357,-216.5,-352,-216.5</points>
<connection>
<GID>233</GID>
<name>OUT_0</name></connection>
<intersection>-352 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-352,-212,-347.5,-212</points>
<connection>
<GID>230</GID>
<name>IN_1</name></connection>
<intersection>-352 0</intersection></hsegment></shape></wire>
<wire>
<ID>104</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-341.5,-211,-336.5,-211</points>
<connection>
<GID>234</GID>
<name>N_in0</name></connection>
<connection>
<GID>230</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>105</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-338.5,-220.5,-338.5,-220</points>
<intersection>-220.5 2</intersection>
<intersection>-220 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-338.5,-220,-336.5,-220</points>
<connection>
<GID>235</GID>
<name>N_in0</name></connection>
<intersection>-338.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-341,-220.5,-338.5,-220.5</points>
<connection>
<GID>231</GID>
<name>OUT</name></connection>
<intersection>-338.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>106</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-352.5,-215.5,-352.5,-210</points>
<intersection>-215.5 3</intersection>
<intersection>-214.5 1</intersection>
<intersection>-210 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-357.5,-214.5,-352.5,-214.5</points>
<connection>
<GID>232</GID>
<name>OUT_0</name></connection>
<intersection>-352.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-352.5,-210,-347.5,-210</points>
<connection>
<GID>230</GID>
<name>IN_0</name></connection>
<intersection>-352.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>-352.5,-215.5,-350.5,-215.5</points>
<connection>
<GID>240</GID>
<name>IN_0</name></connection>
<intersection>-352.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>107</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-346.5,-219.5,-346.5,-215.5</points>
<connection>
<GID>240</GID>
<name>OUT_0</name></connection>
<intersection>-219.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-347,-219.5,-346.5,-219.5</points>
<connection>
<GID>231</GID>
<name>IN_0</name></connection>
<intersection>-346.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>108</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-439.5,-297,-439.5,-283</points>
<intersection>-297 1</intersection>
<intersection>-283 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-439.5,-297,-435,-297</points>
<connection>
<GID>244</GID>
<name>IN_1</name></connection>
<intersection>-439.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-444,-283,-439.5,-283</points>
<connection>
<GID>243</GID>
<name>OUT</name></connection>
<intersection>-439.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>109</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-464,-315.5,-464,-283</points>
<intersection>-315.5 4</intersection>
<intersection>-304 2</intersection>
<intersection>-283 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-464,-283,-463.5,-283</points>
<connection>
<GID>256</GID>
<name>OUT</name></connection>
<intersection>-464 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-464,-304,-434.5,-304</points>
<connection>
<GID>245</GID>
<name>IN_0</name></connection>
<intersection>-464 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-464,-315.5,-436,-315.5</points>
<connection>
<GID>248</GID>
<name>IN_0</name></connection>
<intersection>-464 0</intersection></hsegment></shape></wire>
<wire>
<ID>110</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-453.5,-317.5,-453.5,-279.5</points>
<connection>
<GID>255</GID>
<name>OUT_0</name></connection>
<intersection>-317.5 14</intersection>
<intersection>-306 8</intersection>
<intersection>-283 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-453.5,-283,-450,-283</points>
<intersection>-453.5 0</intersection>
<intersection>-450 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-450,-284,-450,-282</points>
<connection>
<GID>243</GID>
<name>IN_1</name></connection>
<connection>
<GID>243</GID>
<name>IN_0</name></connection>
<intersection>-283 2</intersection></vsegment>
<hsegment>
<ID>8</ID>
<points>-453.5,-306,-434.5,-306</points>
<connection>
<GID>245</GID>
<name>IN_1</name></connection>
<intersection>-453.5 0</intersection></hsegment>
<hsegment>
<ID>14</ID>
<points>-453.5,-317.5,-436,-317.5</points>
<connection>
<GID>248</GID>
<name>IN_1</name></connection>
<intersection>-453.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>111</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-423,-299.5,-423,-296</points>
<intersection>-299.5 1</intersection>
<intersection>-296 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-423,-299.5,-417.5,-299.5</points>
<connection>
<GID>246</GID>
<name>IN_0</name></connection>
<intersection>-423 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-429,-296,-423,-296</points>
<connection>
<GID>244</GID>
<name>OUT</name></connection>
<intersection>-423 0</intersection></hsegment></shape></wire>
<wire>
<ID>112</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-423,-305,-423,-301.5</points>
<intersection>-305 2</intersection>
<intersection>-301.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-423,-301.5,-417.5,-301.5</points>
<connection>
<GID>246</GID>
<name>IN_1</name></connection>
<intersection>-423 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-428.5,-305,-423,-305</points>
<connection>
<GID>245</GID>
<name>OUT</name></connection>
<intersection>-423 0</intersection></hsegment></shape></wire>
<wire>
<ID>113</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-411.5,-300.5,-403.5,-300.5</points>
<connection>
<GID>246</GID>
<name>OUT</name></connection>
<connection>
<GID>247</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>115</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-430,-316.5,-421.5,-316.5</points>
<connection>
<GID>248</GID>
<name>OUT</name></connection>
<intersection>-421.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-421.5,-317.5,-421.5,-315.5</points>
<connection>
<GID>249</GID>
<name>IN_1</name></connection>
<connection>
<GID>249</GID>
<name>IN_0</name></connection>
<intersection>-316.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>116</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-415.5,-316.5,-407,-316.5</points>
<connection>
<GID>249</GID>
<name>OUT</name></connection>
<connection>
<GID>250</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>117</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-472.5,-295,-472.5,-279.5</points>
<connection>
<GID>254</GID>
<name>OUT_0</name></connection>
<intersection>-295 1</intersection>
<intersection>-283 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-472.5,-295,-435,-295</points>
<connection>
<GID>244</GID>
<name>IN_0</name></connection>
<intersection>-472.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-472.5,-283,-469.5,-283</points>
<intersection>-472.5 0</intersection>
<intersection>-469.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-469.5,-284,-469.5,-282</points>
<connection>
<GID>256</GID>
<name>IN_1</name></connection>
<connection>
<GID>256</GID>
<name>IN_0</name></connection>
<intersection>-283 2</intersection></vsegment></shape></wire>
<wire>
<ID>120</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-460.5,-437,-460.5,-383.5</points>
<connection>
<GID>267</GID>
<name>OUT</name></connection>
<intersection>-437 6</intersection>
<intersection>-399.5 4</intersection>
<intersection>-390.5 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>-460.5,-390.5,-402,-390.5</points>
<connection>
<GID>289</GID>
<name>IN_0</name></connection>
<intersection>-460.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-460.5,-399.5,-402,-399.5</points>
<connection>
<GID>291</GID>
<name>IN_0</name></connection>
<intersection>-460.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-460.5,-437,-401.5,-437</points>
<connection>
<GID>299</GID>
<name>IN_0</name></connection>
<intersection>-460.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>121</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-437,-448,-437,-383.5</points>
<intersection>-448 6</intersection>
<intersection>-410 4</intersection>
<intersection>-392.5 2</intersection>
<intersection>-383.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-437,-383.5,-436.5,-383.5</points>
<connection>
<GID>269</GID>
<name>OUT</name></connection>
<intersection>-437 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-437,-392.5,-402,-392.5</points>
<connection>
<GID>289</GID>
<name>IN_1</name></connection>
<intersection>-437 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-437,-410,-402,-410</points>
<connection>
<GID>293</GID>
<name>IN_1</name></connection>
<intersection>-437 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-437,-448,-401.5,-448</points>
<connection>
<GID>297</GID>
<name>IN_1</name></connection>
<intersection>-437 0</intersection></hsegment></shape></wire>
<wire>
<ID>122</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-429.5,-468.5,-429.5,-372.5</points>
<connection>
<GID>265</GID>
<name>OUT_0</name></connection>
<intersection>-468.5 11</intersection>
<intersection>-450 9</intersection>
<intersection>-441 7</intersection>
<intersection>-421 5</intersection>
<intersection>-394.5 1</intersection>
<intersection>-383 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-429.5,-394.5,-402,-394.5</points>
<connection>
<GID>289</GID>
<name>IN_2</name></connection>
<intersection>-429.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-429.5,-383,-421,-383</points>
<intersection>-429.5 0</intersection>
<intersection>-421 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-421,-384,-421,-382</points>
<connection>
<GID>271</GID>
<name>IN_1</name></connection>
<connection>
<GID>271</GID>
<name>IN_0</name></connection>
<intersection>-383 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-429.5,-421,-402,-421</points>
<connection>
<GID>295</GID>
<name>IN_2</name></connection>
<intersection>-429.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-429.5,-441,-401.5,-441</points>
<connection>
<GID>299</GID>
<name>IN_2</name></connection>
<intersection>-429.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-429.5,-450,-401.5,-450</points>
<connection>
<GID>297</GID>
<name>IN_2</name></connection>
<intersection>-429.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-429.5,-468.5,-401.5,-468.5</points>
<connection>
<GID>303</GID>
<name>IN_2</name></connection>
<intersection>-429.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>124</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-450,-466.5,-450,-372.5</points>
<connection>
<GID>263</GID>
<name>OUT_0</name></connection>
<intersection>-466.5 11</intersection>
<intersection>-457 9</intersection>
<intersection>-439 7</intersection>
<intersection>-419 5</intersection>
<intersection>-401.5 1</intersection>
<intersection>-383.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-450,-401.5,-402,-401.5</points>
<connection>
<GID>291</GID>
<name>IN_1</name></connection>
<intersection>-450 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-450,-383.5,-442.5,-383.5</points>
<intersection>-450 0</intersection>
<intersection>-442.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-442.5,-384.5,-442.5,-382.5</points>
<connection>
<GID>269</GID>
<name>IN_1</name></connection>
<connection>
<GID>269</GID>
<name>IN_0</name></connection>
<intersection>-383.5 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-450,-419,-402,-419</points>
<connection>
<GID>295</GID>
<name>IN_1</name></connection>
<intersection>-450 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-450,-439,-401.5,-439</points>
<connection>
<GID>299</GID>
<name>IN_1</name></connection>
<intersection>-450 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-450,-457,-401.5,-457</points>
<connection>
<GID>301</GID>
<name>IN_1</name></connection>
<intersection>-450 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-450,-466.5,-401.5,-466.5</points>
<connection>
<GID>303</GID>
<name>IN_1</name></connection>
<intersection>-450 0</intersection></hsegment></shape></wire>
<wire>
<ID>125</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-414.5,-459,-414.5,-383</points>
<intersection>-459 6</intersection>
<intersection>-412 4</intersection>
<intersection>-403.5 2</intersection>
<intersection>-383 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-415,-383,-414.5,-383</points>
<connection>
<GID>271</GID>
<name>OUT</name></connection>
<intersection>-414.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-414.5,-403.5,-402,-403.5</points>
<connection>
<GID>291</GID>
<name>IN_2</name></connection>
<intersection>-414.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>-414.5,-412,-402,-412</points>
<connection>
<GID>293</GID>
<name>IN_2</name></connection>
<intersection>-414.5 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>-414.5,-459,-401.5,-459</points>
<connection>
<GID>301</GID>
<name>IN_2</name></connection>
<intersection>-414.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>126</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-473.5,-464.5,-473.5,-372.5</points>
<connection>
<GID>261</GID>
<name>OUT_0</name></connection>
<intersection>-464.5 11</intersection>
<intersection>-455 9</intersection>
<intersection>-446 7</intersection>
<intersection>-417 5</intersection>
<intersection>-408 1</intersection>
<intersection>-383.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-473.5,-408,-402,-408</points>
<connection>
<GID>293</GID>
<name>IN_0</name></connection>
<intersection>-473.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-473.5,-383.5,-466.5,-383.5</points>
<intersection>-473.5 0</intersection>
<intersection>-466.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>-466.5,-384.5,-466.5,-382.5</points>
<connection>
<GID>267</GID>
<name>IN_1</name></connection>
<connection>
<GID>267</GID>
<name>IN_0</name></connection>
<intersection>-383.5 2</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>-473.5,-417,-402,-417</points>
<connection>
<GID>295</GID>
<name>IN_0</name></connection>
<intersection>-473.5 0</intersection></hsegment>
<hsegment>
<ID>7</ID>
<points>-473.5,-446,-401.5,-446</points>
<connection>
<GID>297</GID>
<name>IN_0</name></connection>
<intersection>-473.5 0</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>-473.5,-455,-401.5,-455</points>
<connection>
<GID>301</GID>
<name>IN_0</name></connection>
<intersection>-473.5 0</intersection></hsegment>
<hsegment>
<ID>11</ID>
<points>-473.5,-464.5,-401.5,-464.5</points>
<connection>
<GID>303</GID>
<name>IN_0</name></connection>
<intersection>-473.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>131</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-383.5,-401.5,-383.5,-392.5</points>
<intersection>-401.5 1</intersection>
<intersection>-392.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-383.5,-401.5,-364,-401.5</points>
<connection>
<GID>309</GID>
<name>IN_0</name></connection>
<intersection>-383.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-396,-392.5,-383.5,-392.5</points>
<connection>
<GID>289</GID>
<name>OUT</name></connection>
<intersection>-383.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>132</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-383.5,-403.5,-383.5,-401.5</points>
<intersection>-403.5 1</intersection>
<intersection>-401.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-383.5,-403.5,-364,-403.5</points>
<connection>
<GID>309</GID>
<name>IN_1</name></connection>
<intersection>-383.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-396,-401.5,-383.5,-401.5</points>
<connection>
<GID>291</GID>
<name>OUT</name></connection>
<intersection>-383.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>133</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-383.5,-410,-383.5,-405.5</points>
<intersection>-410 2</intersection>
<intersection>-405.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-383.5,-405.5,-364,-405.5</points>
<connection>
<GID>309</GID>
<name>IN_2</name></connection>
<intersection>-383.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-396,-410,-383.5,-410</points>
<connection>
<GID>293</GID>
<name>OUT</name></connection>
<intersection>-383.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>134</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-383.5,-419,-383.5,-407.5</points>
<intersection>-419 2</intersection>
<intersection>-407.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-383.5,-407.5,-364,-407.5</points>
<connection>
<GID>309</GID>
<name>IN_3</name></connection>
<intersection>-383.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-396,-419,-383.5,-419</points>
<connection>
<GID>295</GID>
<name>OUT</name></connection>
<intersection>-383.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>135</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-381,-449.5,-381,-439</points>
<intersection>-449.5 1</intersection>
<intersection>-439 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-381,-449.5,-366.5,-449.5</points>
<connection>
<GID>307</GID>
<name>IN_0</name></connection>
<intersection>-381 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-395.5,-439,-381,-439</points>
<connection>
<GID>299</GID>
<name>OUT</name></connection>
<intersection>-381 0</intersection></hsegment></shape></wire>
<wire>
<ID>136</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-381,-451.5,-381,-448</points>
<intersection>-451.5 1</intersection>
<intersection>-448 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-381,-451.5,-366.5,-451.5</points>
<connection>
<GID>307</GID>
<name>IN_1</name></connection>
<intersection>-381 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-395.5,-448,-381,-448</points>
<connection>
<GID>297</GID>
<name>OUT</name></connection>
<intersection>-381 0</intersection></hsegment></shape></wire>
<wire>
<ID>137</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-381,-457,-381,-453.5</points>
<intersection>-457 2</intersection>
<intersection>-453.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-381,-453.5,-366.5,-453.5</points>
<connection>
<GID>307</GID>
<name>IN_2</name></connection>
<intersection>-381 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-395.5,-457,-381,-457</points>
<connection>
<GID>301</GID>
<name>OUT</name></connection>
<intersection>-381 0</intersection></hsegment></shape></wire>
<wire>
<ID>138</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>-381,-466.5,-381,-455.5</points>
<intersection>-466.5 2</intersection>
<intersection>-455.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>-381,-455.5,-366.5,-455.5</points>
<connection>
<GID>307</GID>
<name>IN_3</name></connection>
<intersection>-381 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>-395.5,-466.5,-381,-466.5</points>
<connection>
<GID>303</GID>
<name>OUT</name></connection>
<intersection>-381 0</intersection></hsegment></shape></wire>
<wire>
<ID>139</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-358,-404.5,-340.5,-404.5</points>
<connection>
<GID>311</GID>
<name>N_in0</name></connection>
<connection>
<GID>309</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>141</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>-360.5,-452.5,-350,-452.5</points>
<connection>
<GID>317</GID>
<name>N_in0</name></connection>
<connection>
<GID>307</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 1>
<page 2>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 2>
<page 3>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 3>
<page 4>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 4>
<page 5>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 5>
<page 6>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 6>
<page 7>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 7>
<page 8>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 8>
<page 9>
<PageViewport>0,0,145.8,-73.7</PageViewport></page 9></circuit>